/* Machine-generated using Migen */
module top(
	input serial_rx,
	output reg serial_tx,
	input clk125_gtp_p,
	input clk125_gtp_n,
	output [14:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash2x_cs_n,
	inout [1:0] spiflash2x_dq,
	input spiflash2x_wp,
	input spiflash2x_hold,
	output sfp_txp,
	output sfp_txn,
	input sfp_rxp,
	input sfp_rxn,
	input sfp_ctl_los,
	input sfp_ctl_mod_present_n,
	output sfp_ctl_rate_select,
	input sfp_ctl_rate_select1,
	output sfp_ctl_tx_disable,
	input sfp_ctl_tx_fault,
	output sfp_ctl_led,
	output user_led,
	inout i2c_scl,
	inout i2c_sda,
	inout dio0_p,
	inout dio0_n,
	inout dio0_p_1,
	inout dio0_n_1,
	inout dio0_p_2,
	inout dio0_n_2,
	inout dio0_p_3,
	inout dio0_n_3,
	inout dio0_p_4,
	inout dio0_n_4,
	inout dio0_p_5,
	inout dio0_n_5,
	inout dio0_p_6,
	inout dio0_n_6,
	inout dio0_p_7,
	inout dio0_n_7,
	inout dio1_p,
	inout dio1_n,
	inout dio1_p_1,
	inout dio1_n_1,
	inout dio1_p_2,
	inout dio1_n_2,
	inout dio1_p_3,
	inout dio1_n_3,
	inout dio1_p_4,
	inout dio1_n_4,
	inout dio1_p_5,
	inout dio1_n_5,
	inout dio1_p_6,
	inout dio1_n_6,
	inout dio1_p_7,
	inout dio1_n_7,
	output urukul2_spi_p_clk,
	inout urukul2_spi_p_mosi,
	inout urukul2_spi_p_miso,
	output [2:0] urukul2_spi_p_cs_n,
	output urukul2_spi_n_clk,
	inout urukul2_spi_n_mosi,
	inout urukul2_spi_n_miso,
	output [2:0] urukul2_spi_n_cs_n,
	output urukul2_dds_reset_sync_in_p,
	output urukul2_dds_reset_sync_in_n,
	inout urukul2_io_update_p,
	inout urukul2_io_update_n,
	inout urukul2_sw0_p,
	inout urukul2_sw0_n,
	inout urukul2_sw1_p,
	inout urukul2_sw1_n,
	inout urukul2_sw2_p,
	inout urukul2_sw2_n,
	inout urukul2_sw3_p,
	inout urukul2_sw3_n,
	output urukul4_spi_p_clk,
	inout urukul4_spi_p_mosi,
	inout urukul4_spi_p_miso,
	output [2:0] urukul4_spi_p_cs_n,
	output urukul4_spi_n_clk,
	inout urukul4_spi_n_mosi,
	inout urukul4_spi_n_miso,
	output [2:0] urukul4_spi_n_cs_n,
	output urukul4_dds_reset_sync_in_p,
	output urukul4_dds_reset_sync_in_n,
	inout urukul4_io_update_p,
	inout urukul4_io_update_n,
	inout urukul4_sw0_p,
	inout urukul4_sw0_n,
	inout urukul4_sw1_p,
	inout urukul4_sw1_n,
	inout urukul4_sw2_p,
	inout urukul4_sw2_n,
	inout urukul4_sw3_p,
	inout urukul4_sw3_n,
	output urukul6_spi_p_clk,
	inout urukul6_spi_p_mosi,
	inout urukul6_spi_p_miso,
	output [2:0] urukul6_spi_p_cs_n,
	output urukul6_spi_n_clk,
	inout urukul6_spi_n_mosi,
	inout urukul6_spi_n_miso,
	output [2:0] urukul6_spi_n_cs_n,
	output urukul6_dds_reset_sync_in_p,
	output urukul6_dds_reset_sync_in_n,
	inout urukul6_io_update_p,
	inout urukul6_io_update_n,
	inout urukul6_sw0_p,
	inout urukul6_sw0_n,
	inout urukul6_sw1_p,
	inout urukul6_sw1_n,
	inout urukul6_sw2_p,
	inout urukul6_sw2_n,
	inout urukul6_sw3_p,
	inout urukul6_sw3_n,
	input sfp_ctl_los_1,
	input sfp_ctl_mod_present_n_1,
	input sfp_ctl_rate_select_1,
	input sfp_ctl_rate_select1_1,
	input sfp_ctl_tx_disable_1,
	input sfp_ctl_tx_fault_1,
	output sfp_ctl_led_1,
	input sfp_ctl_los_2,
	input sfp_ctl_mod_present_n_2,
	input sfp_ctl_rate_select_2,
	input sfp_ctl_rate_select1_2,
	input sfp_ctl_tx_disable_2,
	input sfp_ctl_tx_fault_2,
	output sfp_ctl_led_2,
	input si5324_clkout_fabric_p,
	input si5324_clkout_fabric_n
);

wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_ibus_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_ibus_err;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_dbus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_dbus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_dbus_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_dbus_err;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_interrupt;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_i_adr_o;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_d_adr_o;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_err;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_re = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_re = 1'd0;
reg [29:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full = 30'd0;
wire [17:0] main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_re = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_tmpu_error = 1'd0;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_sram_bus_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_sram_bus_err = 1'd0;
wire [9:0] main_genericstandalone_genericstandalone_genericstandalone_sram_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_sram_we;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w;
reg [13:0] main_genericstandalone_genericstandalone_genericstandalone_interface_adr = 14'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_interface_we = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w = 8'd0;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r = 32'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_err = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_counter = 2'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full = 32'd4367715;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg = 8'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_eop = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data = 8'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx = 32'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg = 8'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount = 4'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_irq;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_status_re;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_status_r;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_status_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full = 2'd0;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_uart_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_eop = 1'd0;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout;
reg [4:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level = 5'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_r;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout;
reg [4:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level = 5'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume = 4'd0;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_r;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr;
wire [8:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop;
wire [7:0] main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data;
wire main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full = 64'd0;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full = 64'd0;
wire [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_r;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_w = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status = 64'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_irq;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_r;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re = 1'd0;
reg [63:0] main_genericstandalone_genericstandalone_genericstandalone_timer0_value = 64'd0;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire main_genericstandalone_genericstandalone_clk125_buf;
wire main_genericstandalone_genericstandalone_clk125_div2;
wire main_genericstandalone_genericstandalone_mmcm_locked;
wire main_genericstandalone_genericstandalone_mmcm_fb;
wire main_genericstandalone_genericstandalone_mmcm_sys;
wire main_genericstandalone_genericstandalone_mmcm_sys4x;
wire main_genericstandalone_genericstandalone_mmcm_sys4x_dqs;
wire main_genericstandalone_genericstandalone_pll_locked;
wire main_genericstandalone_genericstandalone_pll_fb;
wire main_genericstandalone_genericstandalone_pll_clk200;
wire main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg;
wire main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_meta;
wire main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_unbuf;
reg [3:0] main_genericstandalone_genericstandalone_reset_counter = 4'd15;
reg main_genericstandalone_genericstandalone_ic_reset = 1'd1;
reg [1:0] main_genericstandalone_genericstandalone_ddrphy_storage_full = 2'd0;
wire [1:0] main_genericstandalone_genericstandalone_ddrphy_storage;
reg main_genericstandalone_genericstandalone_ddrphy_re = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_w = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_w = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re;
wire main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_r;
reg main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [14:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cs_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata;
reg main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_sd_clk_se;
reg main_genericstandalone_genericstandalone_ddrphy_oe_dqs = 1'd0;
reg [7:0] main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern = 8'd85;
wire main_genericstandalone_genericstandalone_ddrphy_dqs0;
wire main_genericstandalone_genericstandalone_ddrphy_dqs_t0;
wire main_genericstandalone_genericstandalone_ddrphy_dqs1;
wire main_genericstandalone_genericstandalone_ddrphy_dqs_t1;
reg main_genericstandalone_genericstandalone_ddrphy_oe_dq = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t0;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t1;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t2;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t3;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t4;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t5;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t6;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t7;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t8;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t9;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t10;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t11;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t12;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t13;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t14;
wire main_genericstandalone_genericstandalone_ddrphy_dq_o15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15;
wire main_genericstandalone_genericstandalone_ddrphy_dq_t15;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 = 1'd0;
reg main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 = 1'd0;
wire main_genericstandalone_genericstandalone_ddrphy_oe;
reg [3:0] main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en = 4'd0;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte;
wire main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask;
wire main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata;
reg main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_address;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
reg [3:0] main_genericstandalone_genericstandalone_genericstandalone_storage_full = 4'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_re = 1'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status = 32'd0;
reg [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re = 1'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re;
wire main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_r;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_w = 1'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full = 15'd0;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re = 1'd0;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full = 32'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage;
reg main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status = 32'd0;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_en = 1'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_en = 1'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_valid;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cas_n = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_ras_n = 1'd1;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_we_n = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_en = 1'd0;
wire [3:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_en = 1'd0;
wire [31:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_valid;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_bte;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err = 1'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open;
wire [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle = 1'd1;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit;
reg [14:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 = 15'd0;
reg main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_wait;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_done;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count = 3'd4;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_wait;
wire main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_done;
reg [9:0] main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count = 10'd886;
wire [29:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r;
wire [15:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb;
wire main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack;
reg main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we;
reg [2:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti = 3'd0;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_bte = 2'd0;
wire main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_err;
wire [12:0] main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
wire [127:0] main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r;
reg [15:0] main_genericstandalone_genericstandalone_genericstandalone_data_port_we;
reg [127:0] main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w;
reg main_genericstandalone_genericstandalone_genericstandalone_write_from_slave;
reg [1:0] main_genericstandalone_genericstandalone_genericstandalone_adr_offset_r = 2'd0;
wire [12:0] main_genericstandalone_genericstandalone_genericstandalone_tag_port_adr;
wire [19:0] main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_r;
reg main_genericstandalone_genericstandalone_genericstandalone_tag_port_we;
wire [19:0] main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_w;
wire [18:0] main_genericstandalone_genericstandalone_genericstandalone_tag_do_tag;
wire main_genericstandalone_genericstandalone_genericstandalone_tag_do_dirty;
wire [18:0] main_genericstandalone_genericstandalone_genericstandalone_tag_di_tag;
reg main_genericstandalone_genericstandalone_genericstandalone_tag_di_dirty;
reg main_genericstandalone_genericstandalone_genericstandalone_word_clr;
reg main_genericstandalone_genericstandalone_genericstandalone_word_inc;
reg main_genericstandalone_genericstandalone_clk;
wire [29:0] main_genericstandalone_genericstandalone_spiflash_bus_adr;
wire [31:0] main_genericstandalone_genericstandalone_spiflash_bus_dat_w;
wire [31:0] main_genericstandalone_genericstandalone_spiflash_bus_dat_r;
wire [3:0] main_genericstandalone_genericstandalone_spiflash_bus_sel;
wire main_genericstandalone_genericstandalone_spiflash_bus_cyc;
wire main_genericstandalone_genericstandalone_spiflash_bus_stb;
reg main_genericstandalone_genericstandalone_spiflash_bus_ack = 1'd0;
wire main_genericstandalone_genericstandalone_spiflash_bus_we;
wire [2:0] main_genericstandalone_genericstandalone_spiflash_bus_cti;
wire [1:0] main_genericstandalone_genericstandalone_spiflash_bus_bte;
reg main_genericstandalone_genericstandalone_spiflash_bus_err = 1'd0;
reg [3:0] main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full = 4'd0;
wire [3:0] main_genericstandalone_genericstandalone_spiflash_bitbang_storage;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_re = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_status;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full = 1'd0;
wire main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage;
reg main_genericstandalone_genericstandalone_spiflash_bitbang_en_re = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_cs_n = 1'd1;
reg main_genericstandalone_genericstandalone_spiflash_clk = 1'd0;
reg main_genericstandalone_genericstandalone_spiflash_dq_oe = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_spiflash_o;
reg main_genericstandalone_genericstandalone_spiflash_oe;
wire [1:0] main_genericstandalone_genericstandalone_spiflash_i0;
reg [31:0] main_genericstandalone_genericstandalone_spiflash_sr = 32'd0;
reg main_genericstandalone_genericstandalone_spiflash_i1 = 1'd0;
reg [1:0] main_genericstandalone_genericstandalone_spiflash_dqi = 2'd0;
reg [6:0] main_genericstandalone_genericstandalone_spiflash_counter = 7'd0;
wire main_genericstandalone_genericstandalone_qpll_reset;
wire main_genericstandalone_genericstandalone_qpll_lock;
wire main_genericstandalone_genericstandalone_qpll_clk;
wire main_genericstandalone_genericstandalone_qpll_refclk;
reg main_genericstandalone_pcs_transmitpath_config_stb;
wire [15:0] main_genericstandalone_pcs_transmitpath_config_reg;
wire main_genericstandalone_pcs_transmitpath_tx_stb;
reg main_genericstandalone_pcs_transmitpath_tx_ack;
wire [7:0] main_genericstandalone_pcs_transmitpath_tx_data;
reg [7:0] main_genericstandalone_pcs_transmitpath_d0;
reg main_genericstandalone_pcs_transmitpath_k0;
reg [9:0] main_genericstandalone_pcs_transmitpath_output0 = 10'd0;
reg main_genericstandalone_pcs_transmitpath_disparity = 1'd0;
wire [7:0] main_genericstandalone_pcs_transmitpath_d1;
wire main_genericstandalone_pcs_transmitpath_k1;
reg main_genericstandalone_pcs_transmitpath_disp_in = 1'd0;
reg [9:0] main_genericstandalone_pcs_transmitpath_output1;
reg main_genericstandalone_pcs_transmitpath_disp_out;
reg [5:0] main_genericstandalone_pcs_transmitpath_code6b = 6'd0;
reg main_genericstandalone_pcs_transmitpath_code6b_unbalanced = 1'd0;
reg main_genericstandalone_pcs_transmitpath_code6b_flip = 1'd0;
reg [3:0] main_genericstandalone_pcs_transmitpath_code4b = 4'd0;
reg main_genericstandalone_pcs_transmitpath_code4b_unbalanced = 1'd0;
reg main_genericstandalone_pcs_transmitpath_code4b_flip = 1'd0;
reg main_genericstandalone_pcs_transmitpath_alt7_rd0 = 1'd0;
reg main_genericstandalone_pcs_transmitpath_alt7_rd1 = 1'd0;
reg [5:0] main_genericstandalone_pcs_transmitpath_output_6b;
wire main_genericstandalone_pcs_transmitpath_disp_inter;
reg [3:0] main_genericstandalone_pcs_transmitpath_output_4b;
wire [9:0] main_genericstandalone_pcs_transmitpath_output_msb_first;
reg main_genericstandalone_pcs_transmitpath_parity = 1'd0;
reg main_genericstandalone_pcs_transmitpath_c_type = 1'd0;
reg [15:0] main_genericstandalone_pcs_transmitpath_config_reg_buffer = 16'd0;
reg main_genericstandalone_pcs_transmitpath_load_config_reg_buffer;
reg main_genericstandalone_pcs_receivepath_rx_en;
wire [7:0] main_genericstandalone_pcs_receivepath_rx_data;
reg main_genericstandalone_pcs_receivepath_seen_valid_ci;
reg main_genericstandalone_pcs_receivepath_seen_config_reg = 1'd0;
reg [15:0] main_genericstandalone_pcs_receivepath_config_reg = 16'd0;
wire [9:0] main_genericstandalone_pcs_receivepath_input;
wire [7:0] main_genericstandalone_pcs_receivepath_d;
reg main_genericstandalone_pcs_receivepath_k = 1'd0;
reg [9:0] main_genericstandalone_pcs_receivepath_input_msb_first;
reg [4:0] main_genericstandalone_pcs_receivepath_code5b = 5'd0;
reg [2:0] main_genericstandalone_pcs_receivepath_code3b = 3'd0;
reg [7:0] main_genericstandalone_pcs_receivepath_config_reg_lsb = 8'd0;
reg main_genericstandalone_pcs_receivepath_load_config_reg_lsb;
reg main_genericstandalone_pcs_receivepath_load_config_reg_msb;
reg main_genericstandalone_pcs_receivepath_first_preamble_byte;
wire main_genericstandalone_pcs_sink_stb;
wire main_genericstandalone_pcs_sink_ack;
wire main_genericstandalone_pcs_sink_eop;
wire [7:0] main_genericstandalone_pcs_sink_payload_data;
wire main_genericstandalone_pcs_sink_payload_last_be;
wire main_genericstandalone_pcs_sink_payload_error;
reg main_genericstandalone_pcs_source_stb = 1'd0;
wire main_genericstandalone_pcs_source_ack;
wire main_genericstandalone_pcs_source_eop;
reg [7:0] main_genericstandalone_pcs_source_payload_data = 8'd0;
reg main_genericstandalone_pcs_source_payload_last_be = 1'd0;
reg main_genericstandalone_pcs_source_payload_error = 1'd0;
reg main_genericstandalone_pcs_link_up;
reg main_genericstandalone_pcs_restart;
reg main_genericstandalone_pcs_rx_en_d = 1'd0;
wire main_genericstandalone_pcs_seen_valid_ci_i;
wire main_genericstandalone_pcs_seen_valid_ci_o;
reg main_genericstandalone_pcs_seen_valid_ci_toggle_i = 1'd0;
wire main_genericstandalone_pcs_seen_valid_ci_toggle_o;
reg main_genericstandalone_pcs_seen_valid_ci_toggle_o_r = 1'd0;
reg [19:0] main_genericstandalone_pcs_checker_counter = 20'd0;
reg main_genericstandalone_pcs_checker_tick = 1'd0;
reg main_genericstandalone_pcs_checker_ok = 1'd0;
reg main_genericstandalone_pcs_autoneg_ack;
reg main_genericstandalone_pcs_rx_config_reg_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_o;
reg main_genericstandalone_pcs_rx_config_reg_toggle_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_toggle_o;
reg main_genericstandalone_pcs_rx_config_reg_toggle_o_r = 1'd0;
reg main_genericstandalone_pcs_rx_config_reg_ack_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_ack_o;
reg main_genericstandalone_pcs_rx_config_reg_ack_toggle_i = 1'd0;
wire main_genericstandalone_pcs_rx_config_reg_ack_toggle_o;
reg main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r = 1'd0;
reg main_genericstandalone_pcs_wait;
wire main_genericstandalone_pcs_done;
reg [20:0] main_genericstandalone_pcs_count = 21'd1250000;
reg [2:0] main_genericstandalone_pcs_c_counter = 3'd0;
reg [15:0] main_genericstandalone_pcs_previous_config_reg = 16'd0;
wire eth_tx_clk;
wire eth_tx_rst;
wire eth_rx_clk;
wire eth_rx_rst;
wire eth_tx_half_clk;
wire eth_rx_half_clk;
wire main_genericstandalone_txoutclk;
wire main_genericstandalone_rxoutclk;
wire main_genericstandalone_tx_reset;
wire main_genericstandalone_tx_mmcm_locked;
wire [19:0] main_genericstandalone_tx_data0;
wire main_genericstandalone_tx_reset_done;
wire main_genericstandalone_rx_reset;
wire main_genericstandalone_rx_mmcm_locked;
wire [19:0] main_genericstandalone_rx_data0;
wire main_genericstandalone_rx_reset_done;
wire main_genericstandalone_rx_pma_reset_done;
wire [8:0] main_genericstandalone_drpaddr;
wire main_genericstandalone_drpen;
wire [15:0] main_genericstandalone_drpdi;
wire main_genericstandalone_drprdy;
wire [15:0] main_genericstandalone_drpdo;
wire main_genericstandalone_drpwe;
wire main_genericstandalone_txoutclk_rebuffer;
wire main_genericstandalone_rxoutclk_rebuffer;
wire main_genericstandalone_tx_mmcm_fb;
(* dont_touch = "true" *) reg main_genericstandalone_tx_mmcm_reset = 1'd1;
wire main_genericstandalone_clk_tx_unbuf;
wire main_genericstandalone_clk_tx_half_unbuf;
wire main_genericstandalone_rx_mmcm_fb;
(* dont_touch = "true" *) reg main_genericstandalone_rx_mmcm_reset = 1'd1;
wire main_genericstandalone_clk_rx_unbuf;
wire main_genericstandalone_clk_rx_half_unbuf;
(* dont_touch = "true" *) reg main_genericstandalone_tx_init_qpll_reset0 = 1'd0;
wire main_genericstandalone_tx_init_qpll_lock0;
(* dont_touch = "true" *) reg main_genericstandalone_tx_init_tx_reset0 = 1'd0;
reg main_genericstandalone_tx_init_done;
reg main_genericstandalone_tx_init_qpll_reset1;
reg main_genericstandalone_tx_init_tx_reset1;
wire main_genericstandalone_tx_init_qpll_lock1;
reg [5:0] main_genericstandalone_tx_init_timer = 6'd0;
reg main_genericstandalone_tx_init_tick = 1'd0;
(* dont_touch = "true" *) reg main_genericstandalone_rx_init_rx_reset0 = 1'd0;
wire main_genericstandalone_rx_init_rx_pma_reset_done0;
wire [8:0] main_genericstandalone_rx_init_drpaddr;
reg main_genericstandalone_rx_init_drpen;
reg [15:0] main_genericstandalone_rx_init_drpdi;
wire main_genericstandalone_rx_init_drprdy;
wire [15:0] main_genericstandalone_rx_init_drpdo;
reg main_genericstandalone_rx_init_drpwe;
wire main_genericstandalone_rx_init_enable;
wire main_genericstandalone_rx_init_restart;
reg main_genericstandalone_rx_init_done;
reg main_genericstandalone_rx_init_rx_reset1;
wire main_genericstandalone_rx_init_rx_pma_reset_done1;
reg [15:0] main_genericstandalone_rx_init_drpvalue = 16'd0;
reg main_genericstandalone_rx_init_drpmask;
reg main_genericstandalone_rx_init_rx_pma_reset_done_r = 1'd0;
wire main_genericstandalone_i;
wire main_genericstandalone_o;
reg main_genericstandalone_toggle_i = 1'd0;
wire main_genericstandalone_toggle_o;
reg main_genericstandalone_toggle_o_r = 1'd0;
reg [12:0] main_genericstandalone_cdr_lock_counter = 13'd0;
reg main_genericstandalone_cdr_locked = 1'd0;
wire [9:0] main_genericstandalone_tx_data1;
reg [19:0] main_genericstandalone_tx_data_half = 20'd0;
wire [19:0] main_genericstandalone_rx_data_half;
reg [9:0] main_genericstandalone_rx_data1 = 10'd0;
reg [19:0] main_genericstandalone_buf = 20'd0;
reg main_genericstandalone_phase_half = 1'd0;
reg main_genericstandalone_phase_half_rereg = 1'd0;
wire main_genericstandalone_tx_gap_inserter_sink_stb;
reg main_genericstandalone_tx_gap_inserter_sink_ack;
wire main_genericstandalone_tx_gap_inserter_sink_eop;
wire [7:0] main_genericstandalone_tx_gap_inserter_sink_payload_data;
wire main_genericstandalone_tx_gap_inserter_sink_payload_last_be;
wire main_genericstandalone_tx_gap_inserter_sink_payload_error;
reg main_genericstandalone_tx_gap_inserter_source_stb;
wire main_genericstandalone_tx_gap_inserter_source_ack;
reg main_genericstandalone_tx_gap_inserter_source_eop;
reg [7:0] main_genericstandalone_tx_gap_inserter_source_payload_data;
reg main_genericstandalone_tx_gap_inserter_source_payload_last_be;
reg main_genericstandalone_tx_gap_inserter_source_payload_error;
reg [3:0] main_genericstandalone_tx_gap_inserter_counter = 4'd0;
reg main_genericstandalone_tx_gap_inserter_counter_reset;
reg main_genericstandalone_tx_gap_inserter_counter_ce;
reg [31:0] main_genericstandalone_preamble_errors_status = 32'd0;
reg [31:0] main_genericstandalone_crc_errors_status = 32'd0;
wire main_genericstandalone_preamble_inserter_sink_stb;
reg main_genericstandalone_preamble_inserter_sink_ack;
wire main_genericstandalone_preamble_inserter_sink_eop;
wire [7:0] main_genericstandalone_preamble_inserter_sink_payload_data;
wire main_genericstandalone_preamble_inserter_sink_payload_last_be;
wire main_genericstandalone_preamble_inserter_sink_payload_error;
reg main_genericstandalone_preamble_inserter_source_stb;
wire main_genericstandalone_preamble_inserter_source_ack;
reg main_genericstandalone_preamble_inserter_source_eop;
reg [7:0] main_genericstandalone_preamble_inserter_source_payload_data;
wire main_genericstandalone_preamble_inserter_source_payload_last_be;
reg main_genericstandalone_preamble_inserter_source_payload_error;
reg [63:0] main_genericstandalone_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] main_genericstandalone_preamble_inserter_cnt = 3'd0;
reg main_genericstandalone_preamble_inserter_clr_cnt;
reg main_genericstandalone_preamble_inserter_inc_cnt;
wire main_genericstandalone_preamble_checker_sink_stb;
reg main_genericstandalone_preamble_checker_sink_ack;
wire main_genericstandalone_preamble_checker_sink_eop;
wire [7:0] main_genericstandalone_preamble_checker_sink_payload_data;
wire main_genericstandalone_preamble_checker_sink_payload_last_be;
wire main_genericstandalone_preamble_checker_sink_payload_error;
reg main_genericstandalone_preamble_checker_source_stb;
wire main_genericstandalone_preamble_checker_source_ack;
reg main_genericstandalone_preamble_checker_source_eop;
wire [7:0] main_genericstandalone_preamble_checker_source_payload_data;
wire main_genericstandalone_preamble_checker_source_payload_last_be;
reg main_genericstandalone_preamble_checker_source_payload_error;
reg main_genericstandalone_preamble_checker_error;
wire main_genericstandalone_crc32_inserter_sink_stb;
reg main_genericstandalone_crc32_inserter_sink_ack;
wire main_genericstandalone_crc32_inserter_sink_eop;
wire [7:0] main_genericstandalone_crc32_inserter_sink_payload_data;
wire main_genericstandalone_crc32_inserter_sink_payload_last_be;
wire main_genericstandalone_crc32_inserter_sink_payload_error;
reg main_genericstandalone_crc32_inserter_source_stb;
wire main_genericstandalone_crc32_inserter_source_ack;
reg main_genericstandalone_crc32_inserter_source_eop;
reg [7:0] main_genericstandalone_crc32_inserter_source_payload_data;
reg main_genericstandalone_crc32_inserter_source_payload_last_be;
reg main_genericstandalone_crc32_inserter_source_payload_error;
reg [7:0] main_genericstandalone_crc32_inserter_data0;
wire [31:0] main_genericstandalone_crc32_inserter_value;
wire main_genericstandalone_crc32_inserter_error;
wire [7:0] main_genericstandalone_crc32_inserter_data1;
wire [31:0] main_genericstandalone_crc32_inserter_last;
reg [31:0] main_genericstandalone_crc32_inserter_next;
reg [31:0] main_genericstandalone_crc32_inserter_reg = 32'd4294967295;
reg main_genericstandalone_crc32_inserter_ce;
reg main_genericstandalone_crc32_inserter_reset;
reg [1:0] main_genericstandalone_crc32_inserter_cnt = 2'd3;
wire main_genericstandalone_crc32_inserter_cnt_done;
reg main_genericstandalone_crc32_inserter_is_ongoing0;
reg main_genericstandalone_crc32_inserter_is_ongoing1;
wire main_genericstandalone_crc32_checker_sink_sink_stb;
reg main_genericstandalone_crc32_checker_sink_sink_ack;
wire main_genericstandalone_crc32_checker_sink_sink_eop;
wire [7:0] main_genericstandalone_crc32_checker_sink_sink_payload_data;
wire main_genericstandalone_crc32_checker_sink_sink_payload_last_be;
wire main_genericstandalone_crc32_checker_sink_sink_payload_error;
wire main_genericstandalone_crc32_checker_source_source_stb;
wire main_genericstandalone_crc32_checker_source_source_ack;
wire main_genericstandalone_crc32_checker_source_source_eop;
wire [7:0] main_genericstandalone_crc32_checker_source_source_payload_data;
wire main_genericstandalone_crc32_checker_source_source_payload_last_be;
reg main_genericstandalone_crc32_checker_source_source_payload_error;
wire main_genericstandalone_crc32_checker_error;
wire [7:0] main_genericstandalone_crc32_checker_crc_data0;
wire [31:0] main_genericstandalone_crc32_checker_crc_value;
wire main_genericstandalone_crc32_checker_crc_error;
wire [7:0] main_genericstandalone_crc32_checker_crc_data1;
wire [31:0] main_genericstandalone_crc32_checker_crc_last;
reg [31:0] main_genericstandalone_crc32_checker_crc_next;
reg [31:0] main_genericstandalone_crc32_checker_crc_reg = 32'd4294967295;
reg main_genericstandalone_crc32_checker_crc_ce;
reg main_genericstandalone_crc32_checker_crc_reset;
reg main_genericstandalone_crc32_checker_syncfifo_sink_stb;
wire main_genericstandalone_crc32_checker_syncfifo_sink_ack;
wire main_genericstandalone_crc32_checker_syncfifo_sink_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_sink_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_sink_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_source_stb;
wire main_genericstandalone_crc32_checker_syncfifo_source_ack;
wire main_genericstandalone_crc32_checker_syncfifo_source_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_source_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_source_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_we;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_re;
wire main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_syncfifo_din;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_level = 3'd0;
reg main_genericstandalone_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] main_genericstandalone_crc32_checker_syncfifo_wrport_adr;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_wrport_dat_r;
wire main_genericstandalone_crc32_checker_syncfifo_wrport_we;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w;
wire main_genericstandalone_crc32_checker_syncfifo_do_read;
wire [2:0] main_genericstandalone_crc32_checker_syncfifo_rdport_adr;
wire [10:0] main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop;
wire [7:0] main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error;
wire main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop;
reg main_genericstandalone_crc32_checker_fifo_reset;
wire main_genericstandalone_crc32_checker_fifo_in;
wire main_genericstandalone_crc32_checker_fifo_out;
wire main_genericstandalone_crc32_checker_fifo_full;
wire main_genericstandalone_ps_preamble_error_i;
wire main_genericstandalone_ps_preamble_error_o;
reg main_genericstandalone_ps_preamble_error_toggle_i = 1'd0;
wire main_genericstandalone_ps_preamble_error_toggle_o;
reg main_genericstandalone_ps_preamble_error_toggle_o_r = 1'd0;
wire main_genericstandalone_ps_crc_error_i;
wire main_genericstandalone_ps_crc_error_o;
reg main_genericstandalone_ps_crc_error_toggle_i = 1'd0;
wire main_genericstandalone_ps_crc_error_toggle_o;
reg main_genericstandalone_ps_crc_error_toggle_o_r = 1'd0;
wire main_genericstandalone_padding_inserter_sink_stb;
reg main_genericstandalone_padding_inserter_sink_ack;
wire main_genericstandalone_padding_inserter_sink_eop;
wire [7:0] main_genericstandalone_padding_inserter_sink_payload_data;
wire main_genericstandalone_padding_inserter_sink_payload_last_be;
wire main_genericstandalone_padding_inserter_sink_payload_error;
reg main_genericstandalone_padding_inserter_source_stb;
wire main_genericstandalone_padding_inserter_source_ack;
reg main_genericstandalone_padding_inserter_source_eop;
reg [7:0] main_genericstandalone_padding_inserter_source_payload_data;
reg main_genericstandalone_padding_inserter_source_payload_last_be;
reg main_genericstandalone_padding_inserter_source_payload_error;
reg [15:0] main_genericstandalone_padding_inserter_counter = 16'd1;
wire main_genericstandalone_padding_inserter_counter_done;
reg main_genericstandalone_padding_inserter_counter_reset;
reg main_genericstandalone_padding_inserter_counter_ce;
wire main_genericstandalone_padding_checker_sink_stb;
wire main_genericstandalone_padding_checker_sink_ack;
wire main_genericstandalone_padding_checker_sink_eop;
wire [7:0] main_genericstandalone_padding_checker_sink_payload_data;
wire main_genericstandalone_padding_checker_sink_payload_last_be;
wire main_genericstandalone_padding_checker_sink_payload_error;
wire main_genericstandalone_padding_checker_source_stb;
wire main_genericstandalone_padding_checker_source_ack;
wire main_genericstandalone_padding_checker_source_eop;
wire [7:0] main_genericstandalone_padding_checker_source_payload_data;
wire main_genericstandalone_padding_checker_source_payload_last_be;
wire main_genericstandalone_padding_checker_source_payload_error;
wire main_genericstandalone_tx_last_be_sink_stb;
wire main_genericstandalone_tx_last_be_sink_ack;
wire main_genericstandalone_tx_last_be_sink_eop;
wire [7:0] main_genericstandalone_tx_last_be_sink_payload_data;
wire main_genericstandalone_tx_last_be_sink_payload_last_be;
wire main_genericstandalone_tx_last_be_sink_payload_error;
wire main_genericstandalone_tx_last_be_source_stb;
wire main_genericstandalone_tx_last_be_source_ack;
wire main_genericstandalone_tx_last_be_source_eop;
wire [7:0] main_genericstandalone_tx_last_be_source_payload_data;
reg main_genericstandalone_tx_last_be_source_payload_last_be = 1'd0;
reg main_genericstandalone_tx_last_be_source_payload_error = 1'd0;
reg main_genericstandalone_tx_last_be_ongoing = 1'd1;
wire main_genericstandalone_rx_last_be_sink_stb;
wire main_genericstandalone_rx_last_be_sink_ack;
wire main_genericstandalone_rx_last_be_sink_eop;
wire [7:0] main_genericstandalone_rx_last_be_sink_payload_data;
wire main_genericstandalone_rx_last_be_sink_payload_last_be;
wire main_genericstandalone_rx_last_be_sink_payload_error;
wire main_genericstandalone_rx_last_be_source_stb;
wire main_genericstandalone_rx_last_be_source_ack;
wire main_genericstandalone_rx_last_be_source_eop;
wire [7:0] main_genericstandalone_rx_last_be_source_payload_data;
reg main_genericstandalone_rx_last_be_source_payload_last_be;
wire main_genericstandalone_rx_last_be_source_payload_error;
wire main_genericstandalone_tx_converter_sink_sink_stb;
wire main_genericstandalone_tx_converter_sink_sink_ack;
wire main_genericstandalone_tx_converter_sink_sink_eop;
wire [31:0] main_genericstandalone_tx_converter_sink_sink_payload_data;
wire [3:0] main_genericstandalone_tx_converter_sink_sink_payload_last_be;
wire [3:0] main_genericstandalone_tx_converter_sink_sink_payload_error;
wire main_genericstandalone_tx_converter_source_source_stb;
wire main_genericstandalone_tx_converter_source_source_ack;
wire main_genericstandalone_tx_converter_source_source_eop;
wire [7:0] main_genericstandalone_tx_converter_source_source_payload_data;
wire main_genericstandalone_tx_converter_source_source_payload_last_be;
wire main_genericstandalone_tx_converter_source_source_payload_error;
wire main_genericstandalone_tx_converter_converter_sink_stb;
wire main_genericstandalone_tx_converter_converter_sink_ack;
wire main_genericstandalone_tx_converter_converter_sink_eop;
reg [39:0] main_genericstandalone_tx_converter_converter_sink_payload_data;
wire main_genericstandalone_tx_converter_converter_source_stb;
wire main_genericstandalone_tx_converter_converter_source_ack;
wire main_genericstandalone_tx_converter_converter_source_eop;
reg [9:0] main_genericstandalone_tx_converter_converter_source_payload_data;
reg [1:0] main_genericstandalone_tx_converter_converter_mux = 2'd0;
wire main_genericstandalone_tx_converter_converter_last;
wire main_genericstandalone_rx_converter_sink_sink_stb;
wire main_genericstandalone_rx_converter_sink_sink_ack;
wire main_genericstandalone_rx_converter_sink_sink_eop;
wire [7:0] main_genericstandalone_rx_converter_sink_sink_payload_data;
wire main_genericstandalone_rx_converter_sink_sink_payload_last_be;
wire main_genericstandalone_rx_converter_sink_sink_payload_error;
wire main_genericstandalone_rx_converter_source_source_stb;
wire main_genericstandalone_rx_converter_source_source_ack;
wire main_genericstandalone_rx_converter_source_source_eop;
reg [31:0] main_genericstandalone_rx_converter_source_source_payload_data;
reg [3:0] main_genericstandalone_rx_converter_source_source_payload_last_be;
reg [3:0] main_genericstandalone_rx_converter_source_source_payload_error;
wire main_genericstandalone_rx_converter_converter_sink_stb;
wire main_genericstandalone_rx_converter_converter_sink_ack;
wire main_genericstandalone_rx_converter_converter_sink_eop;
wire [9:0] main_genericstandalone_rx_converter_converter_sink_payload_data;
wire main_genericstandalone_rx_converter_converter_source_stb;
wire main_genericstandalone_rx_converter_converter_source_ack;
reg main_genericstandalone_rx_converter_converter_source_eop = 1'd0;
reg [39:0] main_genericstandalone_rx_converter_converter_source_payload_data = 40'd0;
reg [1:0] main_genericstandalone_rx_converter_converter_demux = 2'd0;
wire main_genericstandalone_rx_converter_converter_load_part;
reg main_genericstandalone_rx_converter_converter_strobe_all = 1'd0;
wire main_genericstandalone_tx_cdc_sink_stb;
wire main_genericstandalone_tx_cdc_sink_ack;
wire main_genericstandalone_tx_cdc_sink_eop;
wire [31:0] main_genericstandalone_tx_cdc_sink_payload_data;
wire [3:0] main_genericstandalone_tx_cdc_sink_payload_last_be;
wire [3:0] main_genericstandalone_tx_cdc_sink_payload_error;
wire main_genericstandalone_tx_cdc_source_stb;
wire main_genericstandalone_tx_cdc_source_ack;
wire main_genericstandalone_tx_cdc_source_eop;
wire [31:0] main_genericstandalone_tx_cdc_source_payload_data;
wire [3:0] main_genericstandalone_tx_cdc_source_payload_last_be;
wire [3:0] main_genericstandalone_tx_cdc_source_payload_error;
wire main_genericstandalone_tx_cdc_asyncfifo_we;
wire main_genericstandalone_tx_cdc_asyncfifo_writable;
wire main_genericstandalone_tx_cdc_asyncfifo_re;
wire main_genericstandalone_tx_cdc_asyncfifo_readable;
wire [40:0] main_genericstandalone_tx_cdc_asyncfifo_din;
wire [40:0] main_genericstandalone_tx_cdc_asyncfifo_dout;
wire main_genericstandalone_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_genericstandalone_tx_cdc_graycounter0_q_next;
reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_genericstandalone_tx_cdc_graycounter0_q_next_binary;
wire main_genericstandalone_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_genericstandalone_tx_cdc_graycounter1_q_next;
reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_genericstandalone_tx_cdc_graycounter1_q_next_binary;
wire [6:0] main_genericstandalone_tx_cdc_produce_rdomain;
wire [6:0] main_genericstandalone_tx_cdc_consume_wdomain;
wire [5:0] main_genericstandalone_tx_cdc_wrport_adr;
wire [40:0] main_genericstandalone_tx_cdc_wrport_dat_r;
wire main_genericstandalone_tx_cdc_wrport_we;
wire [40:0] main_genericstandalone_tx_cdc_wrport_dat_w;
wire [5:0] main_genericstandalone_tx_cdc_rdport_adr;
wire [40:0] main_genericstandalone_tx_cdc_rdport_dat_r;
wire [31:0] main_genericstandalone_tx_cdc_fifo_in_payload_data;
wire [3:0] main_genericstandalone_tx_cdc_fifo_in_payload_last_be;
wire [3:0] main_genericstandalone_tx_cdc_fifo_in_payload_error;
wire main_genericstandalone_tx_cdc_fifo_in_eop;
wire [31:0] main_genericstandalone_tx_cdc_fifo_out_payload_data;
wire [3:0] main_genericstandalone_tx_cdc_fifo_out_payload_last_be;
wire [3:0] main_genericstandalone_tx_cdc_fifo_out_payload_error;
wire main_genericstandalone_tx_cdc_fifo_out_eop;
wire main_genericstandalone_rx_cdc_sink_stb;
wire main_genericstandalone_rx_cdc_sink_ack;
wire main_genericstandalone_rx_cdc_sink_eop;
wire [31:0] main_genericstandalone_rx_cdc_sink_payload_data;
wire [3:0] main_genericstandalone_rx_cdc_sink_payload_last_be;
wire [3:0] main_genericstandalone_rx_cdc_sink_payload_error;
wire main_genericstandalone_rx_cdc_source_stb;
wire main_genericstandalone_rx_cdc_source_ack;
wire main_genericstandalone_rx_cdc_source_eop;
wire [31:0] main_genericstandalone_rx_cdc_source_payload_data;
wire [3:0] main_genericstandalone_rx_cdc_source_payload_last_be;
wire [3:0] main_genericstandalone_rx_cdc_source_payload_error;
wire main_genericstandalone_rx_cdc_asyncfifo_we;
wire main_genericstandalone_rx_cdc_asyncfifo_writable;
wire main_genericstandalone_rx_cdc_asyncfifo_re;
wire main_genericstandalone_rx_cdc_asyncfifo_readable;
wire [40:0] main_genericstandalone_rx_cdc_asyncfifo_din;
wire [40:0] main_genericstandalone_rx_cdc_asyncfifo_dout;
wire main_genericstandalone_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_genericstandalone_rx_cdc_graycounter0_q_next;
reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_genericstandalone_rx_cdc_graycounter0_q_next_binary;
wire main_genericstandalone_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_genericstandalone_rx_cdc_graycounter1_q_next;
reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_genericstandalone_rx_cdc_graycounter1_q_next_binary;
wire [6:0] main_genericstandalone_rx_cdc_produce_rdomain;
wire [6:0] main_genericstandalone_rx_cdc_consume_wdomain;
wire [5:0] main_genericstandalone_rx_cdc_wrport_adr;
wire [40:0] main_genericstandalone_rx_cdc_wrport_dat_r;
wire main_genericstandalone_rx_cdc_wrport_we;
wire [40:0] main_genericstandalone_rx_cdc_wrport_dat_w;
wire [5:0] main_genericstandalone_rx_cdc_rdport_adr;
wire [40:0] main_genericstandalone_rx_cdc_rdport_dat_r;
wire [31:0] main_genericstandalone_rx_cdc_fifo_in_payload_data;
wire [3:0] main_genericstandalone_rx_cdc_fifo_in_payload_last_be;
wire [3:0] main_genericstandalone_rx_cdc_fifo_in_payload_error;
wire main_genericstandalone_rx_cdc_fifo_in_eop;
wire [31:0] main_genericstandalone_rx_cdc_fifo_out_payload_data;
wire [3:0] main_genericstandalone_rx_cdc_fifo_out_payload_last_be;
wire [3:0] main_genericstandalone_rx_cdc_fifo_out_payload_error;
wire main_genericstandalone_rx_cdc_fifo_out_eop;
wire main_genericstandalone_sink_stb;
wire main_genericstandalone_sink_ack;
wire main_genericstandalone_sink_eop;
wire [31:0] main_genericstandalone_sink_payload_data;
wire [3:0] main_genericstandalone_sink_payload_last_be;
wire [3:0] main_genericstandalone_sink_payload_error;
wire main_genericstandalone_source_stb;
wire main_genericstandalone_source_ack;
wire main_genericstandalone_source_eop;
wire [31:0] main_genericstandalone_source_payload_data;
wire [3:0] main_genericstandalone_source_payload_last_be;
wire [3:0] main_genericstandalone_source_payload_error;
wire [29:0] main_genericstandalone_bus_adr;
wire [31:0] main_genericstandalone_bus_dat_w;
wire [31:0] main_genericstandalone_bus_dat_r;
wire [3:0] main_genericstandalone_bus_sel;
wire main_genericstandalone_bus_cyc;
wire main_genericstandalone_bus_stb;
wire main_genericstandalone_bus_ack;
wire main_genericstandalone_bus_we;
wire [2:0] main_genericstandalone_bus_cti;
wire [1:0] main_genericstandalone_bus_bte;
wire main_genericstandalone_bus_err;
wire main_genericstandalone_writer_sink_sink_stb;
reg main_genericstandalone_writer_sink_sink_ack = 1'd1;
wire main_genericstandalone_writer_sink_sink_eop;
wire [31:0] main_genericstandalone_writer_sink_sink_payload_data;
wire [3:0] main_genericstandalone_writer_sink_sink_payload_last_be;
wire [3:0] main_genericstandalone_writer_sink_sink_payload_error;
wire [1:0] main_genericstandalone_writer_slot_status;
wire [31:0] main_genericstandalone_writer_length_status;
reg [31:0] main_genericstandalone_writer_errors_status = 32'd0;
wire main_genericstandalone_writer_irq;
wire main_genericstandalone_writer_available_status;
wire main_genericstandalone_writer_available_pending;
wire main_genericstandalone_writer_available_trigger;
reg main_genericstandalone_writer_available_clear;
wire main_genericstandalone_writer_status_re;
wire main_genericstandalone_writer_status_r;
wire main_genericstandalone_writer_status_w;
wire main_genericstandalone_writer_pending_re;
wire main_genericstandalone_writer_pending_r;
wire main_genericstandalone_writer_pending_w;
reg main_genericstandalone_writer_storage_full = 1'd0;
wire main_genericstandalone_writer_storage;
reg main_genericstandalone_writer_re = 1'd0;
reg [2:0] main_genericstandalone_writer_increment;
reg [31:0] main_genericstandalone_writer_counter = 32'd0;
reg main_genericstandalone_writer_counter_reset;
reg main_genericstandalone_writer_counter_ce;
reg [1:0] main_genericstandalone_writer_slot = 2'd0;
reg main_genericstandalone_writer_slot_ce;
reg main_genericstandalone_writer_ongoing;
reg main_genericstandalone_writer_fifo_sink_stb;
wire main_genericstandalone_writer_fifo_sink_ack;
reg main_genericstandalone_writer_fifo_sink_eop = 1'd0;
wire [1:0] main_genericstandalone_writer_fifo_sink_payload_slot;
wire [31:0] main_genericstandalone_writer_fifo_sink_payload_length;
wire main_genericstandalone_writer_fifo_source_stb;
wire main_genericstandalone_writer_fifo_source_ack;
wire main_genericstandalone_writer_fifo_source_eop;
wire [1:0] main_genericstandalone_writer_fifo_source_payload_slot;
wire [31:0] main_genericstandalone_writer_fifo_source_payload_length;
wire main_genericstandalone_writer_fifo_syncfifo_we;
wire main_genericstandalone_writer_fifo_syncfifo_writable;
wire main_genericstandalone_writer_fifo_syncfifo_re;
wire main_genericstandalone_writer_fifo_syncfifo_readable;
wire [34:0] main_genericstandalone_writer_fifo_syncfifo_din;
wire [34:0] main_genericstandalone_writer_fifo_syncfifo_dout;
reg [2:0] main_genericstandalone_writer_fifo_level = 3'd0;
reg main_genericstandalone_writer_fifo_replace = 1'd0;
reg [1:0] main_genericstandalone_writer_fifo_produce = 2'd0;
reg [1:0] main_genericstandalone_writer_fifo_consume = 2'd0;
reg [1:0] main_genericstandalone_writer_fifo_wrport_adr;
wire [34:0] main_genericstandalone_writer_fifo_wrport_dat_r;
wire main_genericstandalone_writer_fifo_wrport_we;
wire [34:0] main_genericstandalone_writer_fifo_wrport_dat_w;
wire main_genericstandalone_writer_fifo_do_read;
wire [1:0] main_genericstandalone_writer_fifo_rdport_adr;
wire [34:0] main_genericstandalone_writer_fifo_rdport_dat_r;
wire [1:0] main_genericstandalone_writer_fifo_fifo_in_payload_slot;
wire [31:0] main_genericstandalone_writer_fifo_fifo_in_payload_length;
wire main_genericstandalone_writer_fifo_fifo_in_eop;
wire [1:0] main_genericstandalone_writer_fifo_fifo_out_payload_slot;
wire [31:0] main_genericstandalone_writer_fifo_fifo_out_payload_length;
wire main_genericstandalone_writer_fifo_fifo_out_eop;
reg [8:0] main_genericstandalone_writer_memory0_adr;
wire [31:0] main_genericstandalone_writer_memory0_dat_r;
reg main_genericstandalone_writer_memory0_we;
reg [31:0] main_genericstandalone_writer_memory0_dat_w;
reg [8:0] main_genericstandalone_writer_memory1_adr;
wire [31:0] main_genericstandalone_writer_memory1_dat_r;
reg main_genericstandalone_writer_memory1_we;
reg [31:0] main_genericstandalone_writer_memory1_dat_w;
reg [8:0] main_genericstandalone_writer_memory2_adr;
wire [31:0] main_genericstandalone_writer_memory2_dat_r;
reg main_genericstandalone_writer_memory2_we;
reg [31:0] main_genericstandalone_writer_memory2_dat_w;
reg [8:0] main_genericstandalone_writer_memory3_adr;
wire [31:0] main_genericstandalone_writer_memory3_dat_r;
reg main_genericstandalone_writer_memory3_we;
reg [31:0] main_genericstandalone_writer_memory3_dat_w;
reg main_genericstandalone_reader_source_source_stb;
wire main_genericstandalone_reader_source_source_ack;
reg main_genericstandalone_reader_source_source_eop;
reg [31:0] main_genericstandalone_reader_source_source_payload_data;
reg [3:0] main_genericstandalone_reader_source_source_payload_last_be;
reg [3:0] main_genericstandalone_reader_source_source_payload_error = 4'd0;
wire main_genericstandalone_reader_start_re;
wire main_genericstandalone_reader_start_r;
reg main_genericstandalone_reader_start_w = 1'd0;
wire main_genericstandalone_reader_ready_status;
reg [1:0] main_genericstandalone_reader_slot_storage_full = 2'd0;
wire [1:0] main_genericstandalone_reader_slot_storage;
reg main_genericstandalone_reader_slot_re = 1'd0;
reg [10:0] main_genericstandalone_reader_length_storage_full = 11'd0;
wire [10:0] main_genericstandalone_reader_length_storage;
reg main_genericstandalone_reader_length_re = 1'd0;
wire main_genericstandalone_reader_irq;
wire main_genericstandalone_reader_done_status;
reg main_genericstandalone_reader_done_pending = 1'd0;
reg main_genericstandalone_reader_done_trigger;
reg main_genericstandalone_reader_done_clear;
wire main_genericstandalone_reader_eventmanager_status_re;
wire main_genericstandalone_reader_eventmanager_status_r;
wire main_genericstandalone_reader_eventmanager_status_w;
wire main_genericstandalone_reader_eventmanager_pending_re;
wire main_genericstandalone_reader_eventmanager_pending_r;
wire main_genericstandalone_reader_eventmanager_pending_w;
reg main_genericstandalone_reader_eventmanager_storage_full = 1'd0;
wire main_genericstandalone_reader_eventmanager_storage;
reg main_genericstandalone_reader_eventmanager_re = 1'd0;
wire main_genericstandalone_reader_fifo_sink_stb;
wire main_genericstandalone_reader_fifo_sink_ack;
reg main_genericstandalone_reader_fifo_sink_eop = 1'd0;
wire [1:0] main_genericstandalone_reader_fifo_sink_payload_slot;
wire [10:0] main_genericstandalone_reader_fifo_sink_payload_length;
wire main_genericstandalone_reader_fifo_source_stb;
reg main_genericstandalone_reader_fifo_source_ack;
wire main_genericstandalone_reader_fifo_source_eop;
wire [1:0] main_genericstandalone_reader_fifo_source_payload_slot;
wire [10:0] main_genericstandalone_reader_fifo_source_payload_length;
wire main_genericstandalone_reader_fifo_syncfifo_we;
wire main_genericstandalone_reader_fifo_syncfifo_writable;
wire main_genericstandalone_reader_fifo_syncfifo_re;
wire main_genericstandalone_reader_fifo_syncfifo_readable;
wire [13:0] main_genericstandalone_reader_fifo_syncfifo_din;
wire [13:0] main_genericstandalone_reader_fifo_syncfifo_dout;
reg [2:0] main_genericstandalone_reader_fifo_level = 3'd0;
reg main_genericstandalone_reader_fifo_replace = 1'd0;
reg [1:0] main_genericstandalone_reader_fifo_produce = 2'd0;
reg [1:0] main_genericstandalone_reader_fifo_consume = 2'd0;
reg [1:0] main_genericstandalone_reader_fifo_wrport_adr;
wire [13:0] main_genericstandalone_reader_fifo_wrport_dat_r;
wire main_genericstandalone_reader_fifo_wrport_we;
wire [13:0] main_genericstandalone_reader_fifo_wrport_dat_w;
wire main_genericstandalone_reader_fifo_do_read;
wire [1:0] main_genericstandalone_reader_fifo_rdport_adr;
wire [13:0] main_genericstandalone_reader_fifo_rdport_dat_r;
wire [1:0] main_genericstandalone_reader_fifo_fifo_in_payload_slot;
wire [10:0] main_genericstandalone_reader_fifo_fifo_in_payload_length;
wire main_genericstandalone_reader_fifo_fifo_in_eop;
wire [1:0] main_genericstandalone_reader_fifo_fifo_out_payload_slot;
wire [10:0] main_genericstandalone_reader_fifo_fifo_out_payload_length;
wire main_genericstandalone_reader_fifo_fifo_out_eop;
reg [10:0] main_genericstandalone_reader_counter = 11'd0;
reg main_genericstandalone_reader_counter_reset;
reg main_genericstandalone_reader_counter_ce;
wire main_genericstandalone_reader_last;
reg main_genericstandalone_reader_last_d = 1'd0;
wire [8:0] main_genericstandalone_reader_memory0_adr;
wire [31:0] main_genericstandalone_reader_memory0_dat_r;
wire [8:0] main_genericstandalone_reader_memory1_adr;
wire [31:0] main_genericstandalone_reader_memory1_dat_r;
wire [8:0] main_genericstandalone_reader_memory2_adr;
wire [31:0] main_genericstandalone_reader_memory2_dat_r;
wire [8:0] main_genericstandalone_reader_memory3_adr;
wire [31:0] main_genericstandalone_reader_memory3_dat_r;
wire main_genericstandalone_ev_irq;
wire [29:0] main_genericstandalone_sram0_bus_adr0;
wire [31:0] main_genericstandalone_sram0_bus_dat_w0;
wire [31:0] main_genericstandalone_sram0_bus_dat_r0;
wire [3:0] main_genericstandalone_sram0_bus_sel0;
wire main_genericstandalone_sram0_bus_cyc0;
wire main_genericstandalone_sram0_bus_stb0;
reg main_genericstandalone_sram0_bus_ack0 = 1'd0;
wire main_genericstandalone_sram0_bus_we0;
wire [2:0] main_genericstandalone_sram0_bus_cti0;
wire [1:0] main_genericstandalone_sram0_bus_bte0;
reg main_genericstandalone_sram0_bus_err0 = 1'd0;
wire [8:0] main_genericstandalone_sram0_adr0;
wire [31:0] main_genericstandalone_sram0_dat_r0;
wire [29:0] main_genericstandalone_sram1_bus_adr0;
wire [31:0] main_genericstandalone_sram1_bus_dat_w0;
wire [31:0] main_genericstandalone_sram1_bus_dat_r0;
wire [3:0] main_genericstandalone_sram1_bus_sel0;
wire main_genericstandalone_sram1_bus_cyc0;
wire main_genericstandalone_sram1_bus_stb0;
reg main_genericstandalone_sram1_bus_ack0 = 1'd0;
wire main_genericstandalone_sram1_bus_we0;
wire [2:0] main_genericstandalone_sram1_bus_cti0;
wire [1:0] main_genericstandalone_sram1_bus_bte0;
reg main_genericstandalone_sram1_bus_err0 = 1'd0;
wire [8:0] main_genericstandalone_sram1_adr0;
wire [31:0] main_genericstandalone_sram1_dat_r0;
wire [29:0] main_genericstandalone_sram2_bus_adr0;
wire [31:0] main_genericstandalone_sram2_bus_dat_w0;
wire [31:0] main_genericstandalone_sram2_bus_dat_r0;
wire [3:0] main_genericstandalone_sram2_bus_sel0;
wire main_genericstandalone_sram2_bus_cyc0;
wire main_genericstandalone_sram2_bus_stb0;
reg main_genericstandalone_sram2_bus_ack0 = 1'd0;
wire main_genericstandalone_sram2_bus_we0;
wire [2:0] main_genericstandalone_sram2_bus_cti0;
wire [1:0] main_genericstandalone_sram2_bus_bte0;
reg main_genericstandalone_sram2_bus_err0 = 1'd0;
wire [8:0] main_genericstandalone_sram2_adr0;
wire [31:0] main_genericstandalone_sram2_dat_r0;
wire [29:0] main_genericstandalone_sram3_bus_adr0;
wire [31:0] main_genericstandalone_sram3_bus_dat_w0;
wire [31:0] main_genericstandalone_sram3_bus_dat_r0;
wire [3:0] main_genericstandalone_sram3_bus_sel0;
wire main_genericstandalone_sram3_bus_cyc0;
wire main_genericstandalone_sram3_bus_stb0;
reg main_genericstandalone_sram3_bus_ack0 = 1'd0;
wire main_genericstandalone_sram3_bus_we0;
wire [2:0] main_genericstandalone_sram3_bus_cti0;
wire [1:0] main_genericstandalone_sram3_bus_bte0;
reg main_genericstandalone_sram3_bus_err0 = 1'd0;
wire [8:0] main_genericstandalone_sram3_adr0;
wire [31:0] main_genericstandalone_sram3_dat_r0;
wire [29:0] main_genericstandalone_sram0_bus_adr1;
wire [31:0] main_genericstandalone_sram0_bus_dat_w1;
wire [31:0] main_genericstandalone_sram0_bus_dat_r1;
wire [3:0] main_genericstandalone_sram0_bus_sel1;
wire main_genericstandalone_sram0_bus_cyc1;
wire main_genericstandalone_sram0_bus_stb1;
reg main_genericstandalone_sram0_bus_ack1 = 1'd0;
wire main_genericstandalone_sram0_bus_we1;
wire [2:0] main_genericstandalone_sram0_bus_cti1;
wire [1:0] main_genericstandalone_sram0_bus_bte1;
reg main_genericstandalone_sram0_bus_err1 = 1'd0;
wire [8:0] main_genericstandalone_sram0_adr1;
wire [31:0] main_genericstandalone_sram0_dat_r1;
reg [3:0] main_genericstandalone_sram0_we;
wire [31:0] main_genericstandalone_sram0_dat_w;
wire [29:0] main_genericstandalone_sram1_bus_adr1;
wire [31:0] main_genericstandalone_sram1_bus_dat_w1;
wire [31:0] main_genericstandalone_sram1_bus_dat_r1;
wire [3:0] main_genericstandalone_sram1_bus_sel1;
wire main_genericstandalone_sram1_bus_cyc1;
wire main_genericstandalone_sram1_bus_stb1;
reg main_genericstandalone_sram1_bus_ack1 = 1'd0;
wire main_genericstandalone_sram1_bus_we1;
wire [2:0] main_genericstandalone_sram1_bus_cti1;
wire [1:0] main_genericstandalone_sram1_bus_bte1;
reg main_genericstandalone_sram1_bus_err1 = 1'd0;
wire [8:0] main_genericstandalone_sram1_adr1;
wire [31:0] main_genericstandalone_sram1_dat_r1;
reg [3:0] main_genericstandalone_sram1_we;
wire [31:0] main_genericstandalone_sram1_dat_w;
wire [29:0] main_genericstandalone_sram2_bus_adr1;
wire [31:0] main_genericstandalone_sram2_bus_dat_w1;
wire [31:0] main_genericstandalone_sram2_bus_dat_r1;
wire [3:0] main_genericstandalone_sram2_bus_sel1;
wire main_genericstandalone_sram2_bus_cyc1;
wire main_genericstandalone_sram2_bus_stb1;
reg main_genericstandalone_sram2_bus_ack1 = 1'd0;
wire main_genericstandalone_sram2_bus_we1;
wire [2:0] main_genericstandalone_sram2_bus_cti1;
wire [1:0] main_genericstandalone_sram2_bus_bte1;
reg main_genericstandalone_sram2_bus_err1 = 1'd0;
wire [8:0] main_genericstandalone_sram2_adr1;
wire [31:0] main_genericstandalone_sram2_dat_r1;
reg [3:0] main_genericstandalone_sram2_we;
wire [31:0] main_genericstandalone_sram2_dat_w;
wire [29:0] main_genericstandalone_sram3_bus_adr1;
wire [31:0] main_genericstandalone_sram3_bus_dat_w1;
wire [31:0] main_genericstandalone_sram3_bus_dat_r1;
wire [3:0] main_genericstandalone_sram3_bus_sel1;
wire main_genericstandalone_sram3_bus_cyc1;
wire main_genericstandalone_sram3_bus_stb1;
reg main_genericstandalone_sram3_bus_ack1 = 1'd0;
wire main_genericstandalone_sram3_bus_we1;
wire [2:0] main_genericstandalone_sram3_bus_cti1;
wire [1:0] main_genericstandalone_sram3_bus_bte1;
reg main_genericstandalone_sram3_bus_err1 = 1'd0;
wire [8:0] main_genericstandalone_sram3_adr1;
wire [31:0] main_genericstandalone_sram3_dat_r1;
reg [3:0] main_genericstandalone_sram3_we;
wire [31:0] main_genericstandalone_sram3_dat_w;
reg [7:0] main_genericstandalone_slave_sel;
reg [7:0] main_genericstandalone_slave_sel_r = 8'd0;
reg main_genericstandalone_kernel_cpu_storage_full = 1'd1;
wire main_genericstandalone_kernel_cpu_storage;
reg main_genericstandalone_kernel_cpu_re = 1'd0;
wire sys_kernel_clk;
wire sys_kernel_rst;
wire [29:0] main_genericstandalone_kernel_cpu_ibus_adr;
wire [31:0] main_genericstandalone_kernel_cpu_ibus_dat_w;
wire [31:0] main_genericstandalone_kernel_cpu_ibus_dat_r;
wire [3:0] main_genericstandalone_kernel_cpu_ibus_sel;
wire main_genericstandalone_kernel_cpu_ibus_cyc;
wire main_genericstandalone_kernel_cpu_ibus_stb;
wire main_genericstandalone_kernel_cpu_ibus_ack;
wire main_genericstandalone_kernel_cpu_ibus_we;
wire [2:0] main_genericstandalone_kernel_cpu_ibus_cti;
wire [1:0] main_genericstandalone_kernel_cpu_ibus_bte;
wire main_genericstandalone_kernel_cpu_ibus_err;
wire [29:0] main_genericstandalone_kernel_cpu_dbus_adr;
wire [31:0] main_genericstandalone_kernel_cpu_dbus_dat_w;
wire [31:0] main_genericstandalone_kernel_cpu_dbus_dat_r;
wire [3:0] main_genericstandalone_kernel_cpu_dbus_sel;
wire main_genericstandalone_kernel_cpu_dbus_cyc;
wire main_genericstandalone_kernel_cpu_dbus_stb;
wire main_genericstandalone_kernel_cpu_dbus_ack;
wire main_genericstandalone_kernel_cpu_dbus_we;
wire [2:0] main_genericstandalone_kernel_cpu_dbus_cti;
wire [1:0] main_genericstandalone_kernel_cpu_dbus_bte;
wire main_genericstandalone_kernel_cpu_dbus_err;
reg [31:0] main_genericstandalone_kernel_cpu_interrupt = 32'd0;
wire [31:0] main_genericstandalone_kernel_cpu_i_adr_o;
wire [31:0] main_genericstandalone_kernel_cpu_d_adr_o;
wire [29:0] main_genericstandalone_kernel_cpu_wb_sdram_adr;
wire [31:0] main_genericstandalone_kernel_cpu_wb_sdram_dat_w;
wire [31:0] main_genericstandalone_kernel_cpu_wb_sdram_dat_r;
wire [3:0] main_genericstandalone_kernel_cpu_wb_sdram_sel;
wire main_genericstandalone_kernel_cpu_wb_sdram_cyc;
wire main_genericstandalone_kernel_cpu_wb_sdram_stb;
wire main_genericstandalone_kernel_cpu_wb_sdram_ack;
wire main_genericstandalone_kernel_cpu_wb_sdram_we;
wire [2:0] main_genericstandalone_kernel_cpu_wb_sdram_cti;
wire [1:0] main_genericstandalone_kernel_cpu_wb_sdram_bte;
wire main_genericstandalone_kernel_cpu_wb_sdram_err;
wire [29:0] main_genericstandalone_mailbox_i1_adr;
wire [31:0] main_genericstandalone_mailbox_i1_dat_w;
reg [31:0] main_genericstandalone_mailbox_i1_dat_r = 32'd0;
wire [3:0] main_genericstandalone_mailbox_i1_sel;
wire main_genericstandalone_mailbox_i1_cyc;
wire main_genericstandalone_mailbox_i1_stb;
reg main_genericstandalone_mailbox_i1_ack = 1'd0;
wire main_genericstandalone_mailbox_i1_we;
wire [2:0] main_genericstandalone_mailbox_i1_cti;
wire [1:0] main_genericstandalone_mailbox_i1_bte;
reg main_genericstandalone_mailbox_i1_err = 1'd0;
wire [29:0] main_genericstandalone_mailbox_i2_adr;
wire [31:0] main_genericstandalone_mailbox_i2_dat_w;
reg [31:0] main_genericstandalone_mailbox_i2_dat_r = 32'd0;
wire [3:0] main_genericstandalone_mailbox_i2_sel;
wire main_genericstandalone_mailbox_i2_cyc;
wire main_genericstandalone_mailbox_i2_stb;
reg main_genericstandalone_mailbox_i2_ack = 1'd0;
wire main_genericstandalone_mailbox_i2_we;
wire [2:0] main_genericstandalone_mailbox_i2_cti;
wire [1:0] main_genericstandalone_mailbox_i2_bte;
reg main_genericstandalone_mailbox_i2_err = 1'd0;
reg [31:0] main_genericstandalone_mailbox0 = 32'd0;
reg [31:0] main_genericstandalone_mailbox1 = 32'd0;
reg [31:0] main_genericstandalone_mailbox2 = 32'd0;
reg [7:0] main_add_identifier_storage_full = 8'd0;
wire [7:0] main_add_identifier_storage;
reg main_add_identifier_re = 1'd0;
wire [7:0] main_add_identifier_status;
wire [5:0] main_add_identifier_adr;
wire [7:0] main_add_identifier_dat_r;
reg main_leds_storage_full = 1'd0;
wire main_leds_storage;
reg main_leds_re = 1'd0;
reg [1:0] main_i2c_status0;
reg [1:0] main_i2c_out_storage_full = 2'd0;
wire [1:0] main_i2c_out_storage;
reg main_i2c_out_re = 1'd0;
reg [1:0] main_i2c_oe_storage_full = 2'd0;
wire [1:0] main_i2c_oe_storage;
reg main_i2c_oe_re = 1'd0;
wire main_i2c_tstriple0_o;
wire main_i2c_tstriple0_oe;
wire main_i2c_tstriple0_i;
wire main_i2c_status1;
wire main_i2c_tstriple1_o;
wire main_i2c_tstriple1_oe;
wire main_i2c_tstriple1_i;
wire main_i2c_status2;
reg [7:0] main_inout_8x0_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x0_serdes_i0;
reg main_inout_8x0_serdes_oe = 1'd0;
wire main_inout_8x0_serdes_pad_i0;
wire main_inout_8x0_serdes_pad_o0;
wire [7:0] main_inout_8x0_serdes_i1;
wire main_inout_8x0_serdes_pad_i1;
wire [7:0] main_inout_8x0_serdes_o1;
wire main_inout_8x0_serdes_t_in;
wire main_inout_8x0_serdes_t_out;
wire main_inout_8x0_serdes_pad_o1;
reg main_inout_8x0_inout_8x0_ointerface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_ointerface0_busy = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_data = 2'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_address = 2'd0;
reg [2:0] main_inout_8x0_inout_8x0_ointerface0_fine_ts = 3'd0;
reg main_inout_8x0_inout_8x0_iinterface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_iinterface0_data = 1'd0;
reg [2:0] main_inout_8x0_inout_8x0_iinterface0_fine_ts = 3'd0;
wire main_inout_8x0_inout_8x0_override_en;
wire main_inout_8x0_inout_8x0_override_o;
wire main_inout_8x0_inout_8x0_override_oe;
wire main_inout_8x0_inout_8x0_input_state;
reg main_inout_8x0_inout_8x0_previous_data = 1'd0;
reg main_inout_8x0_inout_8x0_oe_k = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_sensitivity = 2'd0;
reg main_inout_8x0_inout_8x0_sample = 1'd0;
reg main_inout_8x0_inout_8x0_i_d = 1'd0;
wire [7:0] main_inout_8x0_inout_8x0_i;
reg [2:0] main_inout_8x0_inout_8x0_o;
wire main_inout_8x0_inout_8x0_n;
reg [7:0] main_inout_8x1_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x1_serdes_i0;
reg main_inout_8x1_serdes_oe = 1'd0;
wire main_inout_8x1_serdes_pad_i0;
wire main_inout_8x1_serdes_pad_o0;
wire [7:0] main_inout_8x1_serdes_i1;
wire main_inout_8x1_serdes_pad_i1;
wire [7:0] main_inout_8x1_serdes_o1;
wire main_inout_8x1_serdes_t_in;
wire main_inout_8x1_serdes_t_out;
wire main_inout_8x1_serdes_pad_o1;
reg main_inout_8x1_inout_8x1_ointerface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_ointerface1_busy = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_data = 2'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_address = 2'd0;
reg [2:0] main_inout_8x1_inout_8x1_ointerface1_fine_ts = 3'd0;
reg main_inout_8x1_inout_8x1_iinterface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_iinterface1_data = 1'd0;
reg [2:0] main_inout_8x1_inout_8x1_iinterface1_fine_ts = 3'd0;
wire main_inout_8x1_inout_8x1_override_en;
wire main_inout_8x1_inout_8x1_override_o;
wire main_inout_8x1_inout_8x1_override_oe;
wire main_inout_8x1_inout_8x1_input_state;
reg main_inout_8x1_inout_8x1_previous_data = 1'd0;
reg main_inout_8x1_inout_8x1_oe_k = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_sensitivity = 2'd0;
reg main_inout_8x1_inout_8x1_sample = 1'd0;
reg main_inout_8x1_inout_8x1_i_d = 1'd0;
wire [7:0] main_inout_8x1_inout_8x1_i;
reg [2:0] main_inout_8x1_inout_8x1_o;
wire main_inout_8x1_inout_8x1_n;
reg [7:0] main_inout_8x2_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x2_serdes_i0;
reg main_inout_8x2_serdes_oe = 1'd0;
wire main_inout_8x2_serdes_pad_i0;
wire main_inout_8x2_serdes_pad_o0;
wire [7:0] main_inout_8x2_serdes_i1;
wire main_inout_8x2_serdes_pad_i1;
wire [7:0] main_inout_8x2_serdes_o1;
wire main_inout_8x2_serdes_t_in;
wire main_inout_8x2_serdes_t_out;
wire main_inout_8x2_serdes_pad_o1;
reg main_inout_8x2_inout_8x2_ointerface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_ointerface2_busy = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_data = 2'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_address = 2'd0;
reg [2:0] main_inout_8x2_inout_8x2_ointerface2_fine_ts = 3'd0;
reg main_inout_8x2_inout_8x2_iinterface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_iinterface2_data = 1'd0;
reg [2:0] main_inout_8x2_inout_8x2_iinterface2_fine_ts = 3'd0;
wire main_inout_8x2_inout_8x2_override_en;
wire main_inout_8x2_inout_8x2_override_o;
wire main_inout_8x2_inout_8x2_override_oe;
wire main_inout_8x2_inout_8x2_input_state;
reg main_inout_8x2_inout_8x2_previous_data = 1'd0;
reg main_inout_8x2_inout_8x2_oe_k = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_sensitivity = 2'd0;
reg main_inout_8x2_inout_8x2_sample = 1'd0;
reg main_inout_8x2_inout_8x2_i_d = 1'd0;
wire [7:0] main_inout_8x2_inout_8x2_i;
reg [2:0] main_inout_8x2_inout_8x2_o;
wire main_inout_8x2_inout_8x2_n;
reg [7:0] main_inout_8x3_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x3_serdes_i0;
reg main_inout_8x3_serdes_oe = 1'd0;
wire main_inout_8x3_serdes_pad_i0;
wire main_inout_8x3_serdes_pad_o0;
wire [7:0] main_inout_8x3_serdes_i1;
wire main_inout_8x3_serdes_pad_i1;
wire [7:0] main_inout_8x3_serdes_o1;
wire main_inout_8x3_serdes_t_in;
wire main_inout_8x3_serdes_t_out;
wire main_inout_8x3_serdes_pad_o1;
reg main_inout_8x3_inout_8x3_ointerface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_ointerface3_busy = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_data = 2'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_address = 2'd0;
reg [2:0] main_inout_8x3_inout_8x3_ointerface3_fine_ts = 3'd0;
reg main_inout_8x3_inout_8x3_iinterface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_iinterface3_data = 1'd0;
reg [2:0] main_inout_8x3_inout_8x3_iinterface3_fine_ts = 3'd0;
wire main_inout_8x3_inout_8x3_override_en;
wire main_inout_8x3_inout_8x3_override_o;
wire main_inout_8x3_inout_8x3_override_oe;
wire main_inout_8x3_inout_8x3_input_state;
reg main_inout_8x3_inout_8x3_previous_data = 1'd0;
reg main_inout_8x3_inout_8x3_oe_k = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_sensitivity = 2'd0;
reg main_inout_8x3_inout_8x3_sample = 1'd0;
reg main_inout_8x3_inout_8x3_i_d = 1'd0;
wire [7:0] main_inout_8x3_inout_8x3_i;
reg [2:0] main_inout_8x3_inout_8x3_o;
wire main_inout_8x3_inout_8x3_n;
reg [7:0] main_inout_8x4_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x4_serdes_i0;
reg main_inout_8x4_serdes_oe = 1'd0;
wire main_inout_8x4_serdes_pad_i0;
wire main_inout_8x4_serdes_pad_o0;
wire [7:0] main_inout_8x4_serdes_i1;
wire main_inout_8x4_serdes_pad_i1;
wire [7:0] main_inout_8x4_serdes_o1;
wire main_inout_8x4_serdes_t_in;
wire main_inout_8x4_serdes_t_out;
wire main_inout_8x4_serdes_pad_o1;
reg main_inout_8x4_inout_8x4_ointerface4_stb = 1'd0;
reg main_inout_8x4_inout_8x4_ointerface4_busy = 1'd0;
reg [1:0] main_inout_8x4_inout_8x4_ointerface4_data = 2'd0;
reg [1:0] main_inout_8x4_inout_8x4_ointerface4_address = 2'd0;
reg [2:0] main_inout_8x4_inout_8x4_ointerface4_fine_ts = 3'd0;
reg main_inout_8x4_inout_8x4_iinterface4_stb = 1'd0;
reg main_inout_8x4_inout_8x4_iinterface4_data = 1'd0;
reg [2:0] main_inout_8x4_inout_8x4_iinterface4_fine_ts = 3'd0;
wire main_inout_8x4_inout_8x4_override_en;
wire main_inout_8x4_inout_8x4_override_o;
wire main_inout_8x4_inout_8x4_override_oe;
wire main_inout_8x4_inout_8x4_input_state;
reg main_inout_8x4_inout_8x4_previous_data = 1'd0;
reg main_inout_8x4_inout_8x4_oe_k = 1'd0;
reg [1:0] main_inout_8x4_inout_8x4_sensitivity = 2'd0;
reg main_inout_8x4_inout_8x4_sample = 1'd0;
reg main_inout_8x4_inout_8x4_i_d = 1'd0;
wire [7:0] main_inout_8x4_inout_8x4_i;
reg [2:0] main_inout_8x4_inout_8x4_o;
wire main_inout_8x4_inout_8x4_n;
reg [7:0] main_inout_8x5_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x5_serdes_i0;
reg main_inout_8x5_serdes_oe = 1'd0;
wire main_inout_8x5_serdes_pad_i0;
wire main_inout_8x5_serdes_pad_o0;
wire [7:0] main_inout_8x5_serdes_i1;
wire main_inout_8x5_serdes_pad_i1;
wire [7:0] main_inout_8x5_serdes_o1;
wire main_inout_8x5_serdes_t_in;
wire main_inout_8x5_serdes_t_out;
wire main_inout_8x5_serdes_pad_o1;
reg main_inout_8x5_inout_8x5_ointerface5_stb = 1'd0;
reg main_inout_8x5_inout_8x5_ointerface5_busy = 1'd0;
reg [1:0] main_inout_8x5_inout_8x5_ointerface5_data = 2'd0;
reg [1:0] main_inout_8x5_inout_8x5_ointerface5_address = 2'd0;
reg [2:0] main_inout_8x5_inout_8x5_ointerface5_fine_ts = 3'd0;
reg main_inout_8x5_inout_8x5_iinterface5_stb = 1'd0;
reg main_inout_8x5_inout_8x5_iinterface5_data = 1'd0;
reg [2:0] main_inout_8x5_inout_8x5_iinterface5_fine_ts = 3'd0;
wire main_inout_8x5_inout_8x5_override_en;
wire main_inout_8x5_inout_8x5_override_o;
wire main_inout_8x5_inout_8x5_override_oe;
wire main_inout_8x5_inout_8x5_input_state;
reg main_inout_8x5_inout_8x5_previous_data = 1'd0;
reg main_inout_8x5_inout_8x5_oe_k = 1'd0;
reg [1:0] main_inout_8x5_inout_8x5_sensitivity = 2'd0;
reg main_inout_8x5_inout_8x5_sample = 1'd0;
reg main_inout_8x5_inout_8x5_i_d = 1'd0;
wire [7:0] main_inout_8x5_inout_8x5_i;
reg [2:0] main_inout_8x5_inout_8x5_o;
wire main_inout_8x5_inout_8x5_n;
reg [7:0] main_inout_8x6_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x6_serdes_i0;
reg main_inout_8x6_serdes_oe = 1'd0;
wire main_inout_8x6_serdes_pad_i0;
wire main_inout_8x6_serdes_pad_o0;
wire [7:0] main_inout_8x6_serdes_i1;
wire main_inout_8x6_serdes_pad_i1;
wire [7:0] main_inout_8x6_serdes_o1;
wire main_inout_8x6_serdes_t_in;
wire main_inout_8x6_serdes_t_out;
wire main_inout_8x6_serdes_pad_o1;
reg main_inout_8x6_inout_8x6_ointerface6_stb = 1'd0;
reg main_inout_8x6_inout_8x6_ointerface6_busy = 1'd0;
reg [1:0] main_inout_8x6_inout_8x6_ointerface6_data = 2'd0;
reg [1:0] main_inout_8x6_inout_8x6_ointerface6_address = 2'd0;
reg [2:0] main_inout_8x6_inout_8x6_ointerface6_fine_ts = 3'd0;
reg main_inout_8x6_inout_8x6_iinterface6_stb = 1'd0;
reg main_inout_8x6_inout_8x6_iinterface6_data = 1'd0;
reg [2:0] main_inout_8x6_inout_8x6_iinterface6_fine_ts = 3'd0;
wire main_inout_8x6_inout_8x6_override_en;
wire main_inout_8x6_inout_8x6_override_o;
wire main_inout_8x6_inout_8x6_override_oe;
wire main_inout_8x6_inout_8x6_input_state;
reg main_inout_8x6_inout_8x6_previous_data = 1'd0;
reg main_inout_8x6_inout_8x6_oe_k = 1'd0;
reg [1:0] main_inout_8x6_inout_8x6_sensitivity = 2'd0;
reg main_inout_8x6_inout_8x6_sample = 1'd0;
reg main_inout_8x6_inout_8x6_i_d = 1'd0;
wire [7:0] main_inout_8x6_inout_8x6_i;
reg [2:0] main_inout_8x6_inout_8x6_o;
wire main_inout_8x6_inout_8x6_n;
reg [7:0] main_inout_8x7_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x7_serdes_i0;
reg main_inout_8x7_serdes_oe = 1'd0;
wire main_inout_8x7_serdes_pad_i0;
wire main_inout_8x7_serdes_pad_o0;
wire [7:0] main_inout_8x7_serdes_i1;
wire main_inout_8x7_serdes_pad_i1;
wire [7:0] main_inout_8x7_serdes_o1;
wire main_inout_8x7_serdes_t_in;
wire main_inout_8x7_serdes_t_out;
wire main_inout_8x7_serdes_pad_o1;
reg main_inout_8x7_inout_8x7_ointerface7_stb = 1'd0;
reg main_inout_8x7_inout_8x7_ointerface7_busy = 1'd0;
reg [1:0] main_inout_8x7_inout_8x7_ointerface7_data = 2'd0;
reg [1:0] main_inout_8x7_inout_8x7_ointerface7_address = 2'd0;
reg [2:0] main_inout_8x7_inout_8x7_ointerface7_fine_ts = 3'd0;
reg main_inout_8x7_inout_8x7_iinterface7_stb = 1'd0;
reg main_inout_8x7_inout_8x7_iinterface7_data = 1'd0;
reg [2:0] main_inout_8x7_inout_8x7_iinterface7_fine_ts = 3'd0;
wire main_inout_8x7_inout_8x7_override_en;
wire main_inout_8x7_inout_8x7_override_o;
wire main_inout_8x7_inout_8x7_override_oe;
wire main_inout_8x7_inout_8x7_input_state;
reg main_inout_8x7_inout_8x7_previous_data = 1'd0;
reg main_inout_8x7_inout_8x7_oe_k = 1'd0;
reg [1:0] main_inout_8x7_inout_8x7_sensitivity = 2'd0;
reg main_inout_8x7_inout_8x7_sample = 1'd0;
reg main_inout_8x7_inout_8x7_i_d = 1'd0;
wire [7:0] main_inout_8x7_inout_8x7_i;
reg [2:0] main_inout_8x7_inout_8x7_o;
wire main_inout_8x7_inout_8x7_n;
reg [7:0] main_output_8x0_o = 8'd0;
reg main_output_8x0_t_in = 1'd0;
wire main_output_8x0_t_out;
wire main_output_8x0_pad_o;
reg main_output_8x0_stb = 1'd0;
reg main_output_8x0_busy = 1'd0;
reg main_output_8x0_data = 1'd0;
reg [2:0] main_output_8x0_fine_ts = 3'd0;
wire main_output_8x0_override_en;
wire main_output_8x0_override_o;
reg main_output_8x0_previous_data = 1'd0;
reg [7:0] main_output_8x1_o = 8'd0;
reg main_output_8x1_t_in = 1'd0;
wire main_output_8x1_t_out;
wire main_output_8x1_pad_o;
reg main_output_8x1_stb = 1'd0;
reg main_output_8x1_busy = 1'd0;
reg main_output_8x1_data = 1'd0;
reg [2:0] main_output_8x1_fine_ts = 3'd0;
wire main_output_8x1_override_en;
wire main_output_8x1_override_o;
reg main_output_8x1_previous_data = 1'd0;
reg [7:0] main_output_8x2_o = 8'd0;
reg main_output_8x2_t_in = 1'd0;
wire main_output_8x2_t_out;
wire main_output_8x2_pad_o;
reg main_output_8x2_stb = 1'd0;
reg main_output_8x2_busy = 1'd0;
reg main_output_8x2_data = 1'd0;
reg [2:0] main_output_8x2_fine_ts = 3'd0;
wire main_output_8x2_override_en;
wire main_output_8x2_override_o;
reg main_output_8x2_previous_data = 1'd0;
reg [7:0] main_output_8x3_o = 8'd0;
reg main_output_8x3_t_in = 1'd0;
wire main_output_8x3_t_out;
wire main_output_8x3_pad_o;
reg main_output_8x3_stb = 1'd0;
reg main_output_8x3_busy = 1'd0;
reg main_output_8x3_data = 1'd0;
reg [2:0] main_output_8x3_fine_ts = 3'd0;
wire main_output_8x3_override_en;
wire main_output_8x3_override_o;
reg main_output_8x3_previous_data = 1'd0;
reg [7:0] main_output_8x4_o = 8'd0;
reg main_output_8x4_t_in = 1'd0;
wire main_output_8x4_t_out;
wire main_output_8x4_pad_o;
reg main_output_8x4_stb = 1'd0;
reg main_output_8x4_busy = 1'd0;
reg main_output_8x4_data = 1'd0;
reg [2:0] main_output_8x4_fine_ts = 3'd0;
wire main_output_8x4_override_en;
wire main_output_8x4_override_o;
reg main_output_8x4_previous_data = 1'd0;
reg [7:0] main_output_8x5_o = 8'd0;
reg main_output_8x5_t_in = 1'd0;
wire main_output_8x5_t_out;
wire main_output_8x5_pad_o;
reg main_output_8x5_stb = 1'd0;
reg main_output_8x5_busy = 1'd0;
reg main_output_8x5_data = 1'd0;
reg [2:0] main_output_8x5_fine_ts = 3'd0;
wire main_output_8x5_override_en;
wire main_output_8x5_override_o;
reg main_output_8x5_previous_data = 1'd0;
reg [7:0] main_output_8x6_o = 8'd0;
reg main_output_8x6_t_in = 1'd0;
wire main_output_8x6_t_out;
wire main_output_8x6_pad_o;
reg main_output_8x6_stb = 1'd0;
reg main_output_8x6_busy = 1'd0;
reg main_output_8x6_data = 1'd0;
reg [2:0] main_output_8x6_fine_ts = 3'd0;
wire main_output_8x6_override_en;
wire main_output_8x6_override_o;
reg main_output_8x6_previous_data = 1'd0;
reg [7:0] main_output_8x7_o = 8'd0;
reg main_output_8x7_t_in = 1'd0;
wire main_output_8x7_t_out;
wire main_output_8x7_pad_o;
reg main_output_8x7_stb = 1'd0;
reg main_output_8x7_busy = 1'd0;
reg main_output_8x7_data = 1'd0;
reg [2:0] main_output_8x7_fine_ts = 3'd0;
wire main_output_8x7_override_en;
wire main_output_8x7_override_o;
reg main_output_8x7_previous_data = 1'd0;
wire [2:0] main_spimaster0_interface_cs0;
wire [2:0] main_spimaster0_interface_cs_polarity;
wire main_spimaster0_interface_clk_next;
wire main_spimaster0_interface_clk_polarity;
wire main_spimaster0_interface_cs_next;
wire main_spimaster0_interface_ce;
wire main_spimaster0_interface_sample;
wire main_spimaster0_interface_offline;
wire main_spimaster0_interface_half_duplex;
wire main_spimaster0_interface_sdi;
wire main_spimaster0_interface_sdo;
reg [2:0] main_spimaster0_interface_cs1 = 3'd7;
reg main_spimaster0_interface_clk = 1'd0;
wire main_spimaster0_interface_miso;
wire main_spimaster0_interface_mosi;
reg main_spimaster0_interface_miso_reg = 1'd0;
reg main_spimaster0_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster0_spimachine0_length;
wire main_spimaster0_spimachine0_clk_phase;
reg main_spimaster0_spimachine0_clk_next;
reg main_spimaster0_spimachine0_cs_next;
wire main_spimaster0_spimachine0_ce;
reg main_spimaster0_spimachine0_idle;
wire main_spimaster0_spimachine0_load0;
reg main_spimaster0_spimachine0_readable;
reg main_spimaster0_spimachine0_writable;
wire main_spimaster0_spimachine0_end0;
wire [31:0] main_spimaster0_spimachine0_pdo;
wire [31:0] main_spimaster0_spimachine0_pdi;
reg main_spimaster0_spimachine0_sdo = 1'd0;
wire main_spimaster0_spimachine0_sdi;
wire main_spimaster0_spimachine0_lsb_first;
reg main_spimaster0_spimachine0_load1;
reg main_spimaster0_spimachine0_shift;
reg main_spimaster0_spimachine0_sample;
reg [31:0] main_spimaster0_spimachine0_sr = 32'd0;
wire [7:0] main_spimaster0_spimachine0_div;
reg main_spimaster0_spimachine0_extend;
wire main_spimaster0_spimachine0_done;
reg main_spimaster0_spimachine0_count;
reg [6:0] main_spimaster0_spimachine0_cnt = 7'd0;
wire main_spimaster0_spimachine0_cnt_done;
reg main_spimaster0_spimachine0_do_extend = 1'd0;
reg [4:0] main_spimaster0_spimachine0_n = 5'd0;
reg main_spimaster0_spimachine0_end1 = 1'd0;
reg main_spimaster0_ointerface0_stb = 1'd0;
wire main_spimaster0_ointerface0_busy;
reg [31:0] main_spimaster0_ointerface0_data = 32'd0;
reg main_spimaster0_ointerface0_address = 1'd0;
wire main_spimaster0_iinterface0_stb;
wire [31:0] main_spimaster0_iinterface0_data;
reg main_spimaster0_config_offline = 1'd1;
reg main_spimaster0_config_end = 1'd1;
reg main_spimaster0_config_input = 1'd0;
reg main_spimaster0_config_cs_polarity = 1'd0;
reg main_spimaster0_config_clk_polarity = 1'd0;
reg main_spimaster0_config_clk_phase = 1'd0;
reg main_spimaster0_config_lsb_first = 1'd0;
reg main_spimaster0_config_half_duplex = 1'd0;
reg [4:0] main_spimaster0_config_length = 5'd0;
reg [2:0] main_spimaster0_config_padding = 3'd0;
reg [7:0] main_spimaster0_config_div = 8'd0;
reg [7:0] main_spimaster0_config_cs = 8'd0;
reg main_spimaster0_read = 1'd0;
reg main_pad0 = 1'd0;
reg [7:0] main_output_8x8_o = 8'd0;
reg main_output_8x8_t_in = 1'd0;
wire main_output_8x8_t_out;
wire main_output_8x8_pad_o;
reg main_output_8x8_stb = 1'd0;
reg main_output_8x8_busy = 1'd0;
reg main_output_8x8_data = 1'd0;
reg [2:0] main_output_8x8_fine_ts = 3'd0;
wire main_output_8x8_override_en;
wire main_output_8x8_override_o;
reg main_output_8x8_previous_data = 1'd0;
reg [7:0] main_output_8x9_o = 8'd0;
reg main_output_8x9_t_in = 1'd0;
wire main_output_8x9_t_out;
wire main_output_8x9_pad_o;
reg main_output_8x9_stb = 1'd0;
reg main_output_8x9_busy = 1'd0;
reg main_output_8x9_data = 1'd0;
reg [2:0] main_output_8x9_fine_ts = 3'd0;
wire main_output_8x9_override_en;
wire main_output_8x9_override_o;
reg main_output_8x9_previous_data = 1'd0;
reg [7:0] main_output_8x10_o = 8'd0;
reg main_output_8x10_t_in = 1'd0;
wire main_output_8x10_t_out;
wire main_output_8x10_pad_o;
reg main_output_8x10_stb = 1'd0;
reg main_output_8x10_busy = 1'd0;
reg main_output_8x10_data = 1'd0;
reg [2:0] main_output_8x10_fine_ts = 3'd0;
wire main_output_8x10_override_en;
wire main_output_8x10_override_o;
reg main_output_8x10_previous_data = 1'd0;
reg [7:0] main_output_8x11_o = 8'd0;
reg main_output_8x11_t_in = 1'd0;
wire main_output_8x11_t_out;
wire main_output_8x11_pad_o;
reg main_output_8x11_stb = 1'd0;
reg main_output_8x11_busy = 1'd0;
reg main_output_8x11_data = 1'd0;
reg [2:0] main_output_8x11_fine_ts = 3'd0;
wire main_output_8x11_override_en;
wire main_output_8x11_override_o;
reg main_output_8x11_previous_data = 1'd0;
reg [7:0] main_output_8x12_o = 8'd0;
reg main_output_8x12_t_in = 1'd0;
wire main_output_8x12_t_out;
wire main_output_8x12_pad_o;
reg main_output_8x12_stb = 1'd0;
reg main_output_8x12_busy = 1'd0;
reg main_output_8x12_data = 1'd0;
reg [2:0] main_output_8x12_fine_ts = 3'd0;
wire main_output_8x12_override_en;
wire main_output_8x12_override_o;
reg main_output_8x12_previous_data = 1'd0;
wire [2:0] main_spimaster1_interface_cs0;
wire [2:0] main_spimaster1_interface_cs_polarity;
wire main_spimaster1_interface_clk_next;
wire main_spimaster1_interface_clk_polarity;
wire main_spimaster1_interface_cs_next;
wire main_spimaster1_interface_ce;
wire main_spimaster1_interface_sample;
wire main_spimaster1_interface_offline;
wire main_spimaster1_interface_half_duplex;
wire main_spimaster1_interface_sdi;
wire main_spimaster1_interface_sdo;
reg [2:0] main_spimaster1_interface_cs1 = 3'd7;
reg main_spimaster1_interface_clk = 1'd0;
wire main_spimaster1_interface_miso;
wire main_spimaster1_interface_mosi;
reg main_spimaster1_interface_miso_reg = 1'd0;
reg main_spimaster1_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster1_spimachine1_length;
wire main_spimaster1_spimachine1_clk_phase;
reg main_spimaster1_spimachine1_clk_next;
reg main_spimaster1_spimachine1_cs_next;
wire main_spimaster1_spimachine1_ce;
reg main_spimaster1_spimachine1_idle;
wire main_spimaster1_spimachine1_load0;
reg main_spimaster1_spimachine1_readable;
reg main_spimaster1_spimachine1_writable;
wire main_spimaster1_spimachine1_end0;
wire [31:0] main_spimaster1_spimachine1_pdo;
wire [31:0] main_spimaster1_spimachine1_pdi;
reg main_spimaster1_spimachine1_sdo = 1'd0;
wire main_spimaster1_spimachine1_sdi;
wire main_spimaster1_spimachine1_lsb_first;
reg main_spimaster1_spimachine1_load1;
reg main_spimaster1_spimachine1_shift;
reg main_spimaster1_spimachine1_sample;
reg [31:0] main_spimaster1_spimachine1_sr = 32'd0;
wire [7:0] main_spimaster1_spimachine1_div;
reg main_spimaster1_spimachine1_extend;
wire main_spimaster1_spimachine1_done;
reg main_spimaster1_spimachine1_count;
reg [6:0] main_spimaster1_spimachine1_cnt = 7'd0;
wire main_spimaster1_spimachine1_cnt_done;
reg main_spimaster1_spimachine1_do_extend = 1'd0;
reg [4:0] main_spimaster1_spimachine1_n = 5'd0;
reg main_spimaster1_spimachine1_end1 = 1'd0;
reg main_spimaster1_ointerface1_stb = 1'd0;
wire main_spimaster1_ointerface1_busy;
reg [31:0] main_spimaster1_ointerface1_data = 32'd0;
reg main_spimaster1_ointerface1_address = 1'd0;
wire main_spimaster1_iinterface1_stb;
wire [31:0] main_spimaster1_iinterface1_data;
reg main_spimaster1_config_offline = 1'd1;
reg main_spimaster1_config_end = 1'd1;
reg main_spimaster1_config_input = 1'd0;
reg main_spimaster1_config_cs_polarity = 1'd0;
reg main_spimaster1_config_clk_polarity = 1'd0;
reg main_spimaster1_config_clk_phase = 1'd0;
reg main_spimaster1_config_lsb_first = 1'd0;
reg main_spimaster1_config_half_duplex = 1'd0;
reg [4:0] main_spimaster1_config_length = 5'd0;
reg [2:0] main_spimaster1_config_padding = 3'd0;
reg [7:0] main_spimaster1_config_div = 8'd0;
reg [7:0] main_spimaster1_config_cs = 8'd0;
reg main_spimaster1_read = 1'd0;
reg main_pad1 = 1'd0;
reg [7:0] main_output_8x13_o = 8'd0;
reg main_output_8x13_t_in = 1'd0;
wire main_output_8x13_t_out;
wire main_output_8x13_pad_o;
reg main_output_8x13_stb = 1'd0;
reg main_output_8x13_busy = 1'd0;
reg main_output_8x13_data = 1'd0;
reg [2:0] main_output_8x13_fine_ts = 3'd0;
wire main_output_8x13_override_en;
wire main_output_8x13_override_o;
reg main_output_8x13_previous_data = 1'd0;
reg [7:0] main_output_8x14_o = 8'd0;
reg main_output_8x14_t_in = 1'd0;
wire main_output_8x14_t_out;
wire main_output_8x14_pad_o;
reg main_output_8x14_stb = 1'd0;
reg main_output_8x14_busy = 1'd0;
reg main_output_8x14_data = 1'd0;
reg [2:0] main_output_8x14_fine_ts = 3'd0;
wire main_output_8x14_override_en;
wire main_output_8x14_override_o;
reg main_output_8x14_previous_data = 1'd0;
reg [7:0] main_output_8x15_o = 8'd0;
reg main_output_8x15_t_in = 1'd0;
wire main_output_8x15_t_out;
wire main_output_8x15_pad_o;
reg main_output_8x15_stb = 1'd0;
reg main_output_8x15_busy = 1'd0;
reg main_output_8x15_data = 1'd0;
reg [2:0] main_output_8x15_fine_ts = 3'd0;
wire main_output_8x15_override_en;
wire main_output_8x15_override_o;
reg main_output_8x15_previous_data = 1'd0;
reg [7:0] main_output_8x16_o = 8'd0;
reg main_output_8x16_t_in = 1'd0;
wire main_output_8x16_t_out;
wire main_output_8x16_pad_o;
reg main_output_8x16_stb = 1'd0;
reg main_output_8x16_busy = 1'd0;
reg main_output_8x16_data = 1'd0;
reg [2:0] main_output_8x16_fine_ts = 3'd0;
wire main_output_8x16_override_en;
wire main_output_8x16_override_o;
reg main_output_8x16_previous_data = 1'd0;
reg [7:0] main_output_8x17_o = 8'd0;
reg main_output_8x17_t_in = 1'd0;
wire main_output_8x17_t_out;
wire main_output_8x17_pad_o;
reg main_output_8x17_stb = 1'd0;
reg main_output_8x17_busy = 1'd0;
reg main_output_8x17_data = 1'd0;
reg [2:0] main_output_8x17_fine_ts = 3'd0;
wire main_output_8x17_override_en;
wire main_output_8x17_override_o;
reg main_output_8x17_previous_data = 1'd0;
wire [2:0] main_spimaster2_interface_cs0;
wire [2:0] main_spimaster2_interface_cs_polarity;
wire main_spimaster2_interface_clk_next;
wire main_spimaster2_interface_clk_polarity;
wire main_spimaster2_interface_cs_next;
wire main_spimaster2_interface_ce;
wire main_spimaster2_interface_sample;
wire main_spimaster2_interface_offline;
wire main_spimaster2_interface_half_duplex;
wire main_spimaster2_interface_sdi;
wire main_spimaster2_interface_sdo;
reg [2:0] main_spimaster2_interface_cs1 = 3'd7;
reg main_spimaster2_interface_clk = 1'd0;
wire main_spimaster2_interface_miso;
wire main_spimaster2_interface_mosi;
reg main_spimaster2_interface_miso_reg = 1'd0;
reg main_spimaster2_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster2_spimachine2_length;
wire main_spimaster2_spimachine2_clk_phase;
reg main_spimaster2_spimachine2_clk_next;
reg main_spimaster2_spimachine2_cs_next;
wire main_spimaster2_spimachine2_ce;
reg main_spimaster2_spimachine2_idle;
wire main_spimaster2_spimachine2_load0;
reg main_spimaster2_spimachine2_readable;
reg main_spimaster2_spimachine2_writable;
wire main_spimaster2_spimachine2_end0;
wire [31:0] main_spimaster2_spimachine2_pdo;
wire [31:0] main_spimaster2_spimachine2_pdi;
reg main_spimaster2_spimachine2_sdo = 1'd0;
wire main_spimaster2_spimachine2_sdi;
wire main_spimaster2_spimachine2_lsb_first;
reg main_spimaster2_spimachine2_load1;
reg main_spimaster2_spimachine2_shift;
reg main_spimaster2_spimachine2_sample;
reg [31:0] main_spimaster2_spimachine2_sr = 32'd0;
wire [7:0] main_spimaster2_spimachine2_div;
reg main_spimaster2_spimachine2_extend;
wire main_spimaster2_spimachine2_done;
reg main_spimaster2_spimachine2_count;
reg [6:0] main_spimaster2_spimachine2_cnt = 7'd0;
wire main_spimaster2_spimachine2_cnt_done;
reg main_spimaster2_spimachine2_do_extend = 1'd0;
reg [4:0] main_spimaster2_spimachine2_n = 5'd0;
reg main_spimaster2_spimachine2_end1 = 1'd0;
reg main_spimaster2_ointerface2_stb = 1'd0;
wire main_spimaster2_ointerface2_busy;
reg [31:0] main_spimaster2_ointerface2_data = 32'd0;
reg main_spimaster2_ointerface2_address = 1'd0;
wire main_spimaster2_iinterface2_stb;
wire [31:0] main_spimaster2_iinterface2_data;
reg main_spimaster2_config_offline = 1'd1;
reg main_spimaster2_config_end = 1'd1;
reg main_spimaster2_config_input = 1'd0;
reg main_spimaster2_config_cs_polarity = 1'd0;
reg main_spimaster2_config_clk_polarity = 1'd0;
reg main_spimaster2_config_clk_phase = 1'd0;
reg main_spimaster2_config_lsb_first = 1'd0;
reg main_spimaster2_config_half_duplex = 1'd0;
reg [4:0] main_spimaster2_config_length = 5'd0;
reg [2:0] main_spimaster2_config_padding = 3'd0;
reg [7:0] main_spimaster2_config_div = 8'd0;
reg [7:0] main_spimaster2_config_cs = 8'd0;
reg main_spimaster2_read = 1'd0;
reg main_pad2 = 1'd0;
reg [7:0] main_output_8x18_o = 8'd0;
reg main_output_8x18_t_in = 1'd0;
wire main_output_8x18_t_out;
wire main_output_8x18_pad_o;
reg main_output_8x18_stb = 1'd0;
reg main_output_8x18_busy = 1'd0;
reg main_output_8x18_data = 1'd0;
reg [2:0] main_output_8x18_fine_ts = 3'd0;
wire main_output_8x18_override_en;
wire main_output_8x18_override_o;
reg main_output_8x18_previous_data = 1'd0;
reg [7:0] main_output_8x19_o = 8'd0;
reg main_output_8x19_t_in = 1'd0;
wire main_output_8x19_t_out;
wire main_output_8x19_pad_o;
reg main_output_8x19_stb = 1'd0;
reg main_output_8x19_busy = 1'd0;
reg main_output_8x19_data = 1'd0;
reg [2:0] main_output_8x19_fine_ts = 3'd0;
wire main_output_8x19_override_en;
wire main_output_8x19_override_o;
reg main_output_8x19_previous_data = 1'd0;
reg [7:0] main_output_8x20_o = 8'd0;
reg main_output_8x20_t_in = 1'd0;
wire main_output_8x20_t_out;
wire main_output_8x20_pad_o;
reg main_output_8x20_stb = 1'd0;
reg main_output_8x20_busy = 1'd0;
reg main_output_8x20_data = 1'd0;
reg [2:0] main_output_8x20_fine_ts = 3'd0;
wire main_output_8x20_override_en;
wire main_output_8x20_override_o;
reg main_output_8x20_previous_data = 1'd0;
reg [7:0] main_output_8x21_o = 8'd0;
reg main_output_8x21_t_in = 1'd0;
wire main_output_8x21_t_out;
wire main_output_8x21_pad_o;
reg main_output_8x21_stb = 1'd0;
reg main_output_8x21_busy = 1'd0;
reg main_output_8x21_data = 1'd0;
reg [2:0] main_output_8x21_fine_ts = 3'd0;
wire main_output_8x21_override_en;
wire main_output_8x21_override_o;
reg main_output_8x21_previous_data = 1'd0;
reg [7:0] main_output_8x22_o = 8'd0;
reg main_output_8x22_t_in = 1'd0;
wire main_output_8x22_t_out;
wire main_output_8x22_pad_o;
reg main_output_8x22_stb = 1'd0;
reg main_output_8x22_busy = 1'd0;
reg main_output_8x22_data = 1'd0;
reg [2:0] main_output_8x22_fine_ts = 3'd0;
wire main_output_8x22_override_en;
wire main_output_8x22_override_o;
reg main_output_8x22_previous_data = 1'd0;
reg main_output0_stb = 1'd0;
reg main_output0_busy = 1'd0;
reg main_output0_data = 1'd0;
reg main_output0_pad_o = 1'd0;
wire main_output0_override_en;
wire main_output0_override_o;
reg main_output0_pad_k = 1'd0;
reg main_output1_stb = 1'd0;
reg main_output1_busy = 1'd0;
reg main_output1_data = 1'd0;
reg main_output1_pad_o = 1'd0;
wire main_output1_override_en;
wire main_output1_override_o;
reg main_output1_pad_k = 1'd0;
reg main_stb = 1'd0;
reg main_busy = 1'd0;
reg [31:0] main_data = 32'd0;
reg main_rtio_crg_storage_full = 1'd1;
wire main_rtio_crg_storage;
reg main_rtio_crg_re = 1'd0;
wire main_rtio_crg_pll_locked_status;
wire rtio_clk;
wire rtio_rst;
wire rtiox4_clk;
wire main_rtio_crg_clk_synth_se;
wire main_rtio_crg_pll_locked;
wire main_rtio_crg_rtio_clk;
wire main_rtio_crg_rtiox4_clk;
wire main_rtio_crg_fb_clk;
reg [60:0] main_rtio_tsc_coarse_ts = 61'd0;
wire [63:0] main_rtio_tsc_full_ts;
wire [60:0] main_rtio_tsc_coarse_ts_sys;
wire [63:0] main_rtio_tsc_full_ts_sys;
reg main_rtio_tsc_load = 1'd0;
reg [60:0] main_rtio_tsc_load_value = 61'd0;
wire [60:0] main_rtio_tsc_i;
reg [60:0] main_rtio_tsc_o = 61'd0;
(* dont_touch = "true" *) reg [60:0] main_rtio_tsc_value_gray_rtio = 61'd0;
wire [60:0] main_rtio_tsc_value_gray_sys;
reg [60:0] main_rtio_tsc_value_sys;
reg [1:0] main_rtio_core_cri_cmd;
wire [23:0] main_rtio_core_cri_chan_sel;
wire [63:0] main_rtio_core_cri_o_timestamp;
wire [511:0] main_rtio_core_cri_o_data;
wire [7:0] main_rtio_core_cri_o_address;
wire [2:0] main_rtio_core_cri_o_status;
reg main_rtio_core_cri_o_buffer_space_valid = 1'd0;
reg [15:0] main_rtio_core_cri_o_buffer_space = 16'd0;
wire [63:0] main_rtio_core_cri_i_timeout;
reg [31:0] main_rtio_core_cri_i_data = 32'd0;
reg [63:0] main_rtio_core_cri_i_timestamp = 64'd0;
reg [3:0] main_rtio_core_cri_i_status = 4'd0;
wire main_rtio_core_reset_re;
wire main_rtio_core_reset_r;
reg main_rtio_core_reset_w = 1'd0;
wire main_rtio_core_reset_phy_re;
wire main_rtio_core_reset_phy_r;
reg main_rtio_core_reset_phy_w = 1'd0;
wire main_rtio_core_async_error_re;
wire [2:0] main_rtio_core_async_error_r;
wire [2:0] main_rtio_core_async_error_w;
reg [15:0] main_rtio_core_collision_channel_status = 16'd0;
reg [15:0] main_rtio_core_busy_channel_status = 16'd0;
reg [15:0] main_rtio_core_sequence_error_channel_status = 16'd0;
(* dont_touch = "true" *) reg main_rtio_core_cmd_reset = 1'd1;
(* dont_touch = "true" *) reg main_rtio_core_cmd_reset_phy = 1'd1;
wire rsys_clk;
wire rsys_rst;
wire rio_clk;
wire rio_rst;
wire rio_phy_clk;
wire rio_phy_rst;
reg main_rtio_core_outputs_lanedistributor_sequence_error = 1'd0;
reg [15:0] main_rtio_core_outputs_lanedistributor_sequence_error_channel = 16'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp = 61'd0;
reg main_rtio_core_outputs_lanedistributor_record0_we;
wire main_rtio_core_outputs_lanedistributor_record0_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record0_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record0_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record0_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record0_payload_data;
reg main_rtio_core_outputs_lanedistributor_record1_we;
wire main_rtio_core_outputs_lanedistributor_record1_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record1_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record1_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record1_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record1_payload_data;
reg main_rtio_core_outputs_lanedistributor_record2_we;
wire main_rtio_core_outputs_lanedistributor_record2_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record2_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record2_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record2_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record2_payload_data;
reg main_rtio_core_outputs_lanedistributor_record3_we;
wire main_rtio_core_outputs_lanedistributor_record3_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record3_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record3_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record3_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record3_payload_data;
reg main_rtio_core_outputs_lanedistributor_record4_we;
wire main_rtio_core_outputs_lanedistributor_record4_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record4_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record4_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record4_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record4_payload_data;
reg main_rtio_core_outputs_lanedistributor_record5_we;
wire main_rtio_core_outputs_lanedistributor_record5_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record5_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record5_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record5_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record5_payload_data;
reg main_rtio_core_outputs_lanedistributor_record6_we;
wire main_rtio_core_outputs_lanedistributor_record6_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record6_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record6_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record6_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record6_payload_data;
reg main_rtio_core_outputs_lanedistributor_record7_we;
wire main_rtio_core_outputs_lanedistributor_record7_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record7_seqn;
wire [5:0] main_rtio_core_outputs_lanedistributor_record7_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
wire [1:0] main_rtio_core_outputs_lanedistributor_record7_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record7_payload_data;
wire main_rtio_core_outputs_lanedistributor_o_status_wait;
reg main_rtio_core_outputs_lanedistributor_o_status_underflow = 1'd0;
reg [2:0] main_rtio_core_outputs_lanedistributor_current_lane = 3'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_coarse_timestamp = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 = 61'd0;
reg [11:0] main_rtio_core_outputs_lanedistributor_seqn = 12'd0;
wire [60:0] main_rtio_core_outputs_lanedistributor_coarse_timestamp;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_min_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_last_minus_timestamp = 62'sd0;
wire [2:0] main_rtio_core_outputs_lanedistributor_current_lane_plus_one;
reg main_rtio_core_outputs_lanedistributor_quash = 1'd0;
wire [5:0] main_rtio_core_outputs_lanedistributor_adr;
wire [13:0] main_rtio_core_outputs_lanedistributor_dat_r;
wire signed [13:0] main_rtio_core_outputs_lanedistributor_compensation;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_last;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min;
reg main_rtio_core_outputs_lanedistributor_force_laneB = 1'd0;
reg main_rtio_core_outputs_lanedistributor_use_laneB;
reg [2:0] main_rtio_core_outputs_lanedistributor_use_lanen;
reg main_rtio_core_outputs_lanedistributor_do_write;
reg main_rtio_core_outputs_lanedistributor_do_underflow;
reg main_rtio_core_outputs_lanedistributor_do_sequence_error;
wire [63:0] main_rtio_core_outputs_lanedistributor_compensated_timestamp;
wire main_rtio_core_outputs_lanedistributor_current_lane_writable;
reg main_rtio_core_outputs_lanedistributor_current_lane_writable_r = 1'd1;
wire main_rtio_core_outputs_record0_we;
wire main_rtio_core_outputs_record0_writable;
wire [11:0] main_rtio_core_outputs_record0_seqn0;
wire [5:0] main_rtio_core_outputs_record0_payload_channel0;
wire [63:0] main_rtio_core_outputs_record0_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record0_payload_address0;
wire [31:0] main_rtio_core_outputs_record0_payload_data0;
wire main_rtio_core_outputs_record1_we;
wire main_rtio_core_outputs_record1_writable;
wire [11:0] main_rtio_core_outputs_record1_seqn0;
wire [5:0] main_rtio_core_outputs_record1_payload_channel0;
wire [63:0] main_rtio_core_outputs_record1_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record1_payload_address0;
wire [31:0] main_rtio_core_outputs_record1_payload_data0;
wire main_rtio_core_outputs_record2_we;
wire main_rtio_core_outputs_record2_writable;
wire [11:0] main_rtio_core_outputs_record2_seqn0;
wire [5:0] main_rtio_core_outputs_record2_payload_channel0;
wire [63:0] main_rtio_core_outputs_record2_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record2_payload_address0;
wire [31:0] main_rtio_core_outputs_record2_payload_data0;
wire main_rtio_core_outputs_record3_we;
wire main_rtio_core_outputs_record3_writable;
wire [11:0] main_rtio_core_outputs_record3_seqn0;
wire [5:0] main_rtio_core_outputs_record3_payload_channel0;
wire [63:0] main_rtio_core_outputs_record3_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record3_payload_address0;
wire [31:0] main_rtio_core_outputs_record3_payload_data0;
wire main_rtio_core_outputs_record4_we;
wire main_rtio_core_outputs_record4_writable;
wire [11:0] main_rtio_core_outputs_record4_seqn0;
wire [5:0] main_rtio_core_outputs_record4_payload_channel0;
wire [63:0] main_rtio_core_outputs_record4_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record4_payload_address0;
wire [31:0] main_rtio_core_outputs_record4_payload_data0;
wire main_rtio_core_outputs_record5_we;
wire main_rtio_core_outputs_record5_writable;
wire [11:0] main_rtio_core_outputs_record5_seqn0;
wire [5:0] main_rtio_core_outputs_record5_payload_channel0;
wire [63:0] main_rtio_core_outputs_record5_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record5_payload_address0;
wire [31:0] main_rtio_core_outputs_record5_payload_data0;
wire main_rtio_core_outputs_record6_we;
wire main_rtio_core_outputs_record6_writable;
wire [11:0] main_rtio_core_outputs_record6_seqn0;
wire [5:0] main_rtio_core_outputs_record6_payload_channel0;
wire [63:0] main_rtio_core_outputs_record6_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record6_payload_address0;
wire [31:0] main_rtio_core_outputs_record6_payload_data0;
wire main_rtio_core_outputs_record7_we;
wire main_rtio_core_outputs_record7_writable;
wire [11:0] main_rtio_core_outputs_record7_seqn0;
wire [5:0] main_rtio_core_outputs_record7_payload_channel0;
wire [63:0] main_rtio_core_outputs_record7_payload_timestamp0;
wire [1:0] main_rtio_core_outputs_record7_payload_address0;
wire [31:0] main_rtio_core_outputs_record7_payload_data0;
wire main_rtio_core_outputs_record0_re;
wire main_rtio_core_outputs_record0_readable;
wire [11:0] main_rtio_core_outputs_record0_seqn1;
wire [5:0] main_rtio_core_outputs_record0_payload_channel1;
wire [63:0] main_rtio_core_outputs_record0_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record0_payload_address1;
wire [31:0] main_rtio_core_outputs_record0_payload_data1;
wire main_rtio_core_outputs_record1_re;
wire main_rtio_core_outputs_record1_readable;
wire [11:0] main_rtio_core_outputs_record1_seqn1;
wire [5:0] main_rtio_core_outputs_record1_payload_channel1;
wire [63:0] main_rtio_core_outputs_record1_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record1_payload_address1;
wire [31:0] main_rtio_core_outputs_record1_payload_data1;
wire main_rtio_core_outputs_record2_re;
wire main_rtio_core_outputs_record2_readable;
wire [11:0] main_rtio_core_outputs_record2_seqn1;
wire [5:0] main_rtio_core_outputs_record2_payload_channel1;
wire [63:0] main_rtio_core_outputs_record2_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record2_payload_address1;
wire [31:0] main_rtio_core_outputs_record2_payload_data1;
wire main_rtio_core_outputs_record3_re;
wire main_rtio_core_outputs_record3_readable;
wire [11:0] main_rtio_core_outputs_record3_seqn1;
wire [5:0] main_rtio_core_outputs_record3_payload_channel1;
wire [63:0] main_rtio_core_outputs_record3_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record3_payload_address1;
wire [31:0] main_rtio_core_outputs_record3_payload_data1;
wire main_rtio_core_outputs_record4_re;
wire main_rtio_core_outputs_record4_readable;
wire [11:0] main_rtio_core_outputs_record4_seqn1;
wire [5:0] main_rtio_core_outputs_record4_payload_channel1;
wire [63:0] main_rtio_core_outputs_record4_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record4_payload_address1;
wire [31:0] main_rtio_core_outputs_record4_payload_data1;
wire main_rtio_core_outputs_record5_re;
wire main_rtio_core_outputs_record5_readable;
wire [11:0] main_rtio_core_outputs_record5_seqn1;
wire [5:0] main_rtio_core_outputs_record5_payload_channel1;
wire [63:0] main_rtio_core_outputs_record5_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record5_payload_address1;
wire [31:0] main_rtio_core_outputs_record5_payload_data1;
wire main_rtio_core_outputs_record6_re;
wire main_rtio_core_outputs_record6_readable;
wire [11:0] main_rtio_core_outputs_record6_seqn1;
wire [5:0] main_rtio_core_outputs_record6_payload_channel1;
wire [63:0] main_rtio_core_outputs_record6_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record6_payload_address1;
wire [31:0] main_rtio_core_outputs_record6_payload_data1;
wire main_rtio_core_outputs_record7_re;
wire main_rtio_core_outputs_record7_readable;
wire [11:0] main_rtio_core_outputs_record7_seqn1;
wire [5:0] main_rtio_core_outputs_record7_payload_channel1;
wire [63:0] main_rtio_core_outputs_record7_payload_timestamp1;
wire [1:0] main_rtio_core_outputs_record7_payload_address1;
wire [31:0] main_rtio_core_outputs_record7_payload_data1;
wire main_rtio_core_outputs_asyncfifobuffered0_re;
reg main_rtio_core_outputs_asyncfifobuffered0_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered0_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
wire main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered0_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered1_re;
reg main_rtio_core_outputs_asyncfifobuffered1_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered1_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
wire main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered1_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered2_re;
reg main_rtio_core_outputs_asyncfifobuffered2_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered2_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
wire main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered2_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered3_re;
reg main_rtio_core_outputs_asyncfifobuffered3_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered3_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
wire main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered3_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered4_re;
reg main_rtio_core_outputs_asyncfifobuffered4_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered4_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
wire main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered4_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered5_re;
reg main_rtio_core_outputs_asyncfifobuffered5_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered5_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
wire main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered5_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered6_re;
reg main_rtio_core_outputs_asyncfifobuffered6_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered6_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
wire main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered6_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered7_re;
reg main_rtio_core_outputs_asyncfifobuffered7_readable = 1'd0;
reg [115:0] main_rtio_core_outputs_asyncfifobuffered7_dout = 116'd0;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
wire main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered7_wrport_we;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
wire [115:0] main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;
wire main_rtio_core_outputs_gates_record0_re;
wire main_rtio_core_outputs_gates_record0_readable;
wire [11:0] main_rtio_core_outputs_gates_record0_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record0_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record0_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record0_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record0_payload_data0;
wire main_rtio_core_outputs_gates_record1_re;
wire main_rtio_core_outputs_gates_record1_readable;
wire [11:0] main_rtio_core_outputs_gates_record1_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record1_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record1_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record1_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record1_payload_data0;
wire main_rtio_core_outputs_gates_record2_re;
wire main_rtio_core_outputs_gates_record2_readable;
wire [11:0] main_rtio_core_outputs_gates_record2_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record2_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record2_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record2_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record2_payload_data0;
wire main_rtio_core_outputs_gates_record3_re;
wire main_rtio_core_outputs_gates_record3_readable;
wire [11:0] main_rtio_core_outputs_gates_record3_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record3_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record3_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record3_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record3_payload_data0;
wire main_rtio_core_outputs_gates_record4_re;
wire main_rtio_core_outputs_gates_record4_readable;
wire [11:0] main_rtio_core_outputs_gates_record4_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record4_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record4_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record4_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record4_payload_data0;
wire main_rtio_core_outputs_gates_record5_re;
wire main_rtio_core_outputs_gates_record5_readable;
wire [11:0] main_rtio_core_outputs_gates_record5_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record5_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record5_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record5_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record5_payload_data0;
wire main_rtio_core_outputs_gates_record6_re;
wire main_rtio_core_outputs_gates_record6_readable;
wire [11:0] main_rtio_core_outputs_gates_record6_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record6_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record6_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record6_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record6_payload_data0;
wire main_rtio_core_outputs_gates_record7_re;
wire main_rtio_core_outputs_gates_record7_readable;
wire [11:0] main_rtio_core_outputs_gates_record7_seqn0;
wire [5:0] main_rtio_core_outputs_gates_record7_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record7_payload_timestamp;
wire [1:0] main_rtio_core_outputs_gates_record7_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record7_payload_data0;
reg main_rtio_core_outputs_gates_record0_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record0_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record0_replace_occured;
wire main_rtio_core_outputs_gates_record0_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record0_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record0_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record0_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record0_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record1_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record1_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record1_replace_occured;
wire main_rtio_core_outputs_gates_record1_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record1_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record1_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record1_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record1_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record2_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record2_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record2_replace_occured;
wire main_rtio_core_outputs_gates_record2_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record2_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record2_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record2_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record2_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record3_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record3_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record3_replace_occured;
wire main_rtio_core_outputs_gates_record3_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record3_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record3_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record3_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record3_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record4_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record4_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record4_replace_occured;
wire main_rtio_core_outputs_gates_record4_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record4_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record4_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record4_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record4_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record5_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record5_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record5_replace_occured;
wire main_rtio_core_outputs_gates_record5_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record5_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record5_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record5_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record5_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record6_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record6_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record6_replace_occured;
wire main_rtio_core_outputs_gates_record6_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record6_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record6_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record6_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record6_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record7_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record7_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record7_replace_occured;
wire main_rtio_core_outputs_gates_record7_nondata_replace_occured;
reg [5:0] main_rtio_core_outputs_gates_record7_payload_channel1 = 6'd0;
reg [2:0] main_rtio_core_outputs_gates_record7_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_gates_record7_payload_address1 = 2'd0;
reg [31:0] main_rtio_core_outputs_gates_record7_payload_data1 = 32'd0;
wire [60:0] main_rtio_core_outputs_gates_coarse_timestamp;
reg main_rtio_core_outputs_collision = 1'd0;
reg [5:0] main_rtio_core_outputs_collision_channel = 6'd0;
reg main_rtio_core_outputs_busy = 1'd0;
reg [5:0] main_rtio_core_outputs_busy_channel = 6'd0;
wire main_rtio_core_outputs_record0_valid0;
wire [11:0] main_rtio_core_outputs_record0_seqn2;
wire main_rtio_core_outputs_record0_replace_occured;
wire main_rtio_core_outputs_record0_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record0_payload_channel2;
wire [2:0] main_rtio_core_outputs_record0_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record0_payload_address2;
wire [31:0] main_rtio_core_outputs_record0_payload_data2;
wire main_rtio_core_outputs_record1_valid0;
wire [11:0] main_rtio_core_outputs_record1_seqn2;
wire main_rtio_core_outputs_record1_replace_occured;
wire main_rtio_core_outputs_record1_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record1_payload_channel2;
wire [2:0] main_rtio_core_outputs_record1_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record1_payload_address2;
wire [31:0] main_rtio_core_outputs_record1_payload_data2;
wire main_rtio_core_outputs_record2_valid0;
wire [11:0] main_rtio_core_outputs_record2_seqn2;
wire main_rtio_core_outputs_record2_replace_occured;
wire main_rtio_core_outputs_record2_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record2_payload_channel2;
wire [2:0] main_rtio_core_outputs_record2_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record2_payload_address2;
wire [31:0] main_rtio_core_outputs_record2_payload_data2;
wire main_rtio_core_outputs_record3_valid0;
wire [11:0] main_rtio_core_outputs_record3_seqn2;
wire main_rtio_core_outputs_record3_replace_occured;
wire main_rtio_core_outputs_record3_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record3_payload_channel2;
wire [2:0] main_rtio_core_outputs_record3_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record3_payload_address2;
wire [31:0] main_rtio_core_outputs_record3_payload_data2;
wire main_rtio_core_outputs_record4_valid0;
wire [11:0] main_rtio_core_outputs_record4_seqn2;
wire main_rtio_core_outputs_record4_replace_occured;
wire main_rtio_core_outputs_record4_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record4_payload_channel2;
wire [2:0] main_rtio_core_outputs_record4_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record4_payload_address2;
wire [31:0] main_rtio_core_outputs_record4_payload_data2;
wire main_rtio_core_outputs_record5_valid0;
wire [11:0] main_rtio_core_outputs_record5_seqn2;
wire main_rtio_core_outputs_record5_replace_occured;
wire main_rtio_core_outputs_record5_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record5_payload_channel2;
wire [2:0] main_rtio_core_outputs_record5_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record5_payload_address2;
wire [31:0] main_rtio_core_outputs_record5_payload_data2;
wire main_rtio_core_outputs_record6_valid0;
wire [11:0] main_rtio_core_outputs_record6_seqn2;
wire main_rtio_core_outputs_record6_replace_occured;
wire main_rtio_core_outputs_record6_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record6_payload_channel2;
wire [2:0] main_rtio_core_outputs_record6_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record6_payload_address2;
wire [31:0] main_rtio_core_outputs_record6_payload_data2;
wire main_rtio_core_outputs_record7_valid0;
wire [11:0] main_rtio_core_outputs_record7_seqn2;
wire main_rtio_core_outputs_record7_replace_occured;
wire main_rtio_core_outputs_record7_nondata_replace_occured;
wire [5:0] main_rtio_core_outputs_record7_payload_channel2;
wire [2:0] main_rtio_core_outputs_record7_payload_fine_ts0;
wire [1:0] main_rtio_core_outputs_record7_payload_address2;
wire [31:0] main_rtio_core_outputs_record7_payload_data2;
reg main_rtio_core_outputs_record0_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record0_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record0_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record0_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record0_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record0_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record0_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record0_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record1_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record1_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record1_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record1_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record1_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record1_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record1_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record1_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record2_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record2_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record2_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record2_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record2_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record2_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record2_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record2_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record3_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record3_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record3_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record3_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record3_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record3_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record3_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record3_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record4_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record4_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record4_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record4_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record4_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record4_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record4_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record4_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record5_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record5_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record5_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record5_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record5_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record5_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record5_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record5_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record6_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record6_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record6_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record6_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record6_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record6_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record6_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record6_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record7_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record7_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record7_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record7_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record7_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record7_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record7_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record7_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference0;
reg main_rtio_core_outputs_nondata_difference1;
reg main_rtio_core_outputs_nondata_difference2;
reg main_rtio_core_outputs_nondata_difference3;
reg main_rtio_core_outputs_record8_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record8_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record8_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record8_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record8_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record8_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record8_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record8_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record9_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record9_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record9_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record9_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record9_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record9_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record9_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record9_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record10_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record10_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record10_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record10_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record10_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record10_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record10_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record10_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record11_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record11_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record11_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record11_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record11_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record11_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record11_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record11_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record12_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record12_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record12_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record12_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record12_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record12_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record12_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record12_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record13_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record13_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record13_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record13_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record13_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record13_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record13_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record13_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record14_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record14_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record14_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record14_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record14_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record14_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record14_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record14_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record15_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record15_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record15_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record15_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record15_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record15_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record15_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record15_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference4;
reg main_rtio_core_outputs_nondata_difference5;
reg main_rtio_core_outputs_nondata_difference6;
reg main_rtio_core_outputs_nondata_difference7;
reg main_rtio_core_outputs_record16_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record16_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record16_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record16_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record16_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record16_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record16_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record16_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record17_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record17_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record17_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record17_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record17_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record17_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record17_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record17_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record18_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record18_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record18_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record18_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record18_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record18_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record18_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record18_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record19_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record19_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record19_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record19_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record19_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record19_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record19_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record19_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record20_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record20_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record20_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record20_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record20_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record20_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record20_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record20_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record21_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record21_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record21_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record21_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record21_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record21_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record21_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record21_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record22_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record22_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record22_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record22_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record22_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record22_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record22_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record22_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record23_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record23_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record23_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record23_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record23_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record23_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record23_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record23_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference8;
reg main_rtio_core_outputs_nondata_difference9;
reg main_rtio_core_outputs_record24_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record24_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record24_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record24_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record24_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record24_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record24_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record24_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record25_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record25_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record25_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record25_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record25_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record25_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record25_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record25_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record26_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record26_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record26_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record26_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record26_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record26_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record26_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record26_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record27_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record27_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record27_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record27_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record27_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record27_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record27_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record27_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record28_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record28_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record28_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record28_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record28_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record28_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record28_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record28_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record29_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record29_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record29_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record29_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record29_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record29_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record29_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record29_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record30_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record30_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record30_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record30_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record30_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record30_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record30_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record30_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record31_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record31_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record31_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record31_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record31_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record31_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record31_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record31_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference10;
reg main_rtio_core_outputs_nondata_difference11;
reg main_rtio_core_outputs_nondata_difference12;
reg main_rtio_core_outputs_nondata_difference13;
reg main_rtio_core_outputs_record32_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record32_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record32_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record32_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record32_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record32_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record32_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record32_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record33_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record33_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record33_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record33_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record33_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record33_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record33_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record33_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record34_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record34_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record34_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record34_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record34_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record34_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record34_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record34_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record35_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record35_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record35_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record35_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record35_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record35_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record35_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record35_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record36_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record36_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record36_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record36_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record36_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record36_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record36_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record36_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record37_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record37_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record37_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record37_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record37_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record37_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record37_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record37_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record38_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record38_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record38_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record38_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record38_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record38_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record38_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record38_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record39_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record39_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record39_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record39_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record39_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record39_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record39_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record39_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference14;
reg main_rtio_core_outputs_nondata_difference15;
reg main_rtio_core_outputs_record40_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record40_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record40_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record40_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record40_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record40_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record40_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record40_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record41_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record41_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record41_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record41_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record41_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record41_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record41_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record41_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record42_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record42_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record42_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record42_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record42_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record42_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record42_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record42_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record43_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record43_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record43_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record43_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record43_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record43_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record43_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record43_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record44_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record44_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record44_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record44_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record44_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record44_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record44_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record44_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record45_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record45_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record45_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record45_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record45_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record45_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record45_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record45_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record46_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record46_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record46_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record46_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record46_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record46_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record46_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record46_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record47_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record47_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record47_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record47_rec_nondata_replace_occured = 1'd0;
reg [5:0] main_rtio_core_outputs_record47_rec_payload_channel = 6'd0;
reg [2:0] main_rtio_core_outputs_record47_rec_payload_fine_ts = 3'd0;
reg [1:0] main_rtio_core_outputs_record47_rec_payload_address = 2'd0;
reg [31:0] main_rtio_core_outputs_record47_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference16;
reg main_rtio_core_outputs_nondata_difference17;
reg main_rtio_core_outputs_nondata_difference18;
reg main_rtio_core_outputs_record0_valid1 = 1'd0;
wire main_rtio_core_outputs_record0_collision;
reg [5:0] main_rtio_core_outputs_record0_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record0_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record0_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record0_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record1_valid1 = 1'd0;
wire main_rtio_core_outputs_record1_collision;
reg [5:0] main_rtio_core_outputs_record1_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record1_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record1_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record1_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record2_valid1 = 1'd0;
wire main_rtio_core_outputs_record2_collision;
reg [5:0] main_rtio_core_outputs_record2_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record2_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record2_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record2_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record3_valid1 = 1'd0;
wire main_rtio_core_outputs_record3_collision;
reg [5:0] main_rtio_core_outputs_record3_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record3_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record3_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record3_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record4_valid1 = 1'd0;
wire main_rtio_core_outputs_record4_collision;
reg [5:0] main_rtio_core_outputs_record4_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record4_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record4_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record4_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record5_valid1 = 1'd0;
wire main_rtio_core_outputs_record5_collision;
reg [5:0] main_rtio_core_outputs_record5_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record5_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record5_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record5_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record6_valid1 = 1'd0;
wire main_rtio_core_outputs_record6_collision;
reg [5:0] main_rtio_core_outputs_record6_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record6_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record6_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record6_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record7_valid1 = 1'd0;
wire main_rtio_core_outputs_record7_collision;
reg [5:0] main_rtio_core_outputs_record7_payload_channel3 = 6'd0;
reg [2:0] main_rtio_core_outputs_record7_payload_fine_ts1 = 3'd0;
reg [1:0] main_rtio_core_outputs_record7_payload_address3 = 2'd0;
reg [31:0] main_rtio_core_outputs_record7_payload_data3 = 32'd0;
reg main_rtio_core_outputs_replace_occured_r0 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r0 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory0_adr;
wire main_rtio_core_outputs_memory0_dat_r;
reg main_rtio_core_outputs_replace_occured_r1 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r1 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory1_adr;
wire main_rtio_core_outputs_memory1_dat_r;
reg main_rtio_core_outputs_replace_occured_r2 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r2 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory2_adr;
wire main_rtio_core_outputs_memory2_dat_r;
reg main_rtio_core_outputs_replace_occured_r3 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r3 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory3_adr;
wire main_rtio_core_outputs_memory3_dat_r;
reg main_rtio_core_outputs_replace_occured_r4 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r4 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory4_adr;
wire main_rtio_core_outputs_memory4_dat_r;
reg main_rtio_core_outputs_replace_occured_r5 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r5 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory5_adr;
wire main_rtio_core_outputs_memory5_dat_r;
reg main_rtio_core_outputs_replace_occured_r6 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r6 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory6_adr;
wire main_rtio_core_outputs_memory6_dat_r;
reg main_rtio_core_outputs_replace_occured_r7 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r7 = 1'd0;
wire [5:0] main_rtio_core_outputs_memory7_adr;
wire main_rtio_core_outputs_memory7_dat_r;
wire main_rtio_core_outputs_selected0;
wire main_rtio_core_outputs_selected1;
wire main_rtio_core_outputs_selected2;
wire main_rtio_core_outputs_selected3;
wire main_rtio_core_outputs_selected4;
wire main_rtio_core_outputs_selected5;
wire main_rtio_core_outputs_selected6;
wire main_rtio_core_outputs_selected7;
wire main_rtio_core_outputs_selected8;
wire main_rtio_core_outputs_selected9;
wire main_rtio_core_outputs_selected10;
wire main_rtio_core_outputs_selected11;
wire main_rtio_core_outputs_selected12;
wire main_rtio_core_outputs_selected13;
wire main_rtio_core_outputs_selected14;
wire main_rtio_core_outputs_selected15;
wire main_rtio_core_outputs_selected16;
wire main_rtio_core_outputs_selected17;
wire main_rtio_core_outputs_selected18;
wire main_rtio_core_outputs_selected19;
wire main_rtio_core_outputs_selected20;
wire main_rtio_core_outputs_selected21;
wire main_rtio_core_outputs_selected22;
wire main_rtio_core_outputs_selected23;
wire main_rtio_core_outputs_selected24;
wire main_rtio_core_outputs_selected25;
wire main_rtio_core_outputs_selected26;
wire main_rtio_core_outputs_selected27;
wire main_rtio_core_outputs_selected28;
wire main_rtio_core_outputs_selected29;
wire main_rtio_core_outputs_selected30;
wire main_rtio_core_outputs_selected31;
wire main_rtio_core_outputs_selected32;
wire main_rtio_core_outputs_selected33;
wire main_rtio_core_outputs_selected34;
wire main_rtio_core_outputs_selected35;
wire main_rtio_core_outputs_selected36;
wire main_rtio_core_outputs_selected37;
wire main_rtio_core_outputs_selected38;
wire main_rtio_core_outputs_selected39;
wire main_rtio_core_outputs_selected40;
wire main_rtio_core_outputs_selected41;
wire main_rtio_core_outputs_selected42;
wire main_rtio_core_outputs_selected43;
wire main_rtio_core_outputs_selected44;
wire main_rtio_core_outputs_selected45;
wire main_rtio_core_outputs_selected46;
wire main_rtio_core_outputs_selected47;
wire main_rtio_core_outputs_selected48;
wire main_rtio_core_outputs_selected49;
wire main_rtio_core_outputs_selected50;
wire main_rtio_core_outputs_selected51;
wire main_rtio_core_outputs_selected52;
wire main_rtio_core_outputs_selected53;
wire main_rtio_core_outputs_selected54;
wire main_rtio_core_outputs_selected55;
wire main_rtio_core_outputs_selected56;
wire main_rtio_core_outputs_selected57;
wire main_rtio_core_outputs_selected58;
wire main_rtio_core_outputs_selected59;
wire main_rtio_core_outputs_selected60;
wire main_rtio_core_outputs_selected61;
wire main_rtio_core_outputs_selected62;
wire main_rtio_core_outputs_selected63;
wire main_rtio_core_outputs_selected64;
wire main_rtio_core_outputs_selected65;
wire main_rtio_core_outputs_selected66;
wire main_rtio_core_outputs_selected67;
wire main_rtio_core_outputs_selected68;
wire main_rtio_core_outputs_selected69;
wire main_rtio_core_outputs_selected70;
wire main_rtio_core_outputs_selected71;
wire main_rtio_core_outputs_selected72;
wire main_rtio_core_outputs_selected73;
wire main_rtio_core_outputs_selected74;
wire main_rtio_core_outputs_selected75;
wire main_rtio_core_outputs_selected76;
wire main_rtio_core_outputs_selected77;
wire main_rtio_core_outputs_selected78;
wire main_rtio_core_outputs_selected79;
wire main_rtio_core_outputs_selected80;
wire main_rtio_core_outputs_selected81;
wire main_rtio_core_outputs_selected82;
wire main_rtio_core_outputs_selected83;
wire main_rtio_core_outputs_selected84;
wire main_rtio_core_outputs_selected85;
wire main_rtio_core_outputs_selected86;
wire main_rtio_core_outputs_selected87;
wire main_rtio_core_outputs_selected88;
wire main_rtio_core_outputs_selected89;
wire main_rtio_core_outputs_selected90;
wire main_rtio_core_outputs_selected91;
wire main_rtio_core_outputs_selected92;
wire main_rtio_core_outputs_selected93;
wire main_rtio_core_outputs_selected94;
wire main_rtio_core_outputs_selected95;
wire main_rtio_core_outputs_selected96;
wire main_rtio_core_outputs_selected97;
wire main_rtio_core_outputs_selected98;
wire main_rtio_core_outputs_selected99;
wire main_rtio_core_outputs_selected100;
wire main_rtio_core_outputs_selected101;
wire main_rtio_core_outputs_selected102;
wire main_rtio_core_outputs_selected103;
wire main_rtio_core_outputs_selected104;
wire main_rtio_core_outputs_selected105;
wire main_rtio_core_outputs_selected106;
wire main_rtio_core_outputs_selected107;
wire main_rtio_core_outputs_selected108;
wire main_rtio_core_outputs_selected109;
wire main_rtio_core_outputs_selected110;
wire main_rtio_core_outputs_selected111;
wire main_rtio_core_outputs_selected112;
wire main_rtio_core_outputs_selected113;
wire main_rtio_core_outputs_selected114;
wire main_rtio_core_outputs_selected115;
wire main_rtio_core_outputs_selected116;
wire main_rtio_core_outputs_selected117;
wire main_rtio_core_outputs_selected118;
wire main_rtio_core_outputs_selected119;
wire main_rtio_core_outputs_selected120;
wire main_rtio_core_outputs_selected121;
wire main_rtio_core_outputs_selected122;
wire main_rtio_core_outputs_selected123;
wire main_rtio_core_outputs_selected124;
wire main_rtio_core_outputs_selected125;
wire main_rtio_core_outputs_selected126;
wire main_rtio_core_outputs_selected127;
wire main_rtio_core_outputs_selected128;
wire main_rtio_core_outputs_selected129;
wire main_rtio_core_outputs_selected130;
wire main_rtio_core_outputs_selected131;
wire main_rtio_core_outputs_selected132;
wire main_rtio_core_outputs_selected133;
wire main_rtio_core_outputs_selected134;
wire main_rtio_core_outputs_selected135;
wire main_rtio_core_outputs_selected136;
wire main_rtio_core_outputs_selected137;
wire main_rtio_core_outputs_selected138;
wire main_rtio_core_outputs_selected139;
wire main_rtio_core_outputs_selected140;
wire main_rtio_core_outputs_selected141;
wire main_rtio_core_outputs_selected142;
wire main_rtio_core_outputs_selected143;
wire main_rtio_core_outputs_selected144;
wire main_rtio_core_outputs_selected145;
wire main_rtio_core_outputs_selected146;
wire main_rtio_core_outputs_selected147;
wire main_rtio_core_outputs_selected148;
wire main_rtio_core_outputs_selected149;
wire main_rtio_core_outputs_selected150;
wire main_rtio_core_outputs_selected151;
wire main_rtio_core_outputs_selected152;
wire main_rtio_core_outputs_selected153;
wire main_rtio_core_outputs_selected154;
wire main_rtio_core_outputs_selected155;
wire main_rtio_core_outputs_selected156;
wire main_rtio_core_outputs_selected157;
wire main_rtio_core_outputs_selected158;
wire main_rtio_core_outputs_selected159;
wire main_rtio_core_outputs_selected160;
wire main_rtio_core_outputs_selected161;
wire main_rtio_core_outputs_selected162;
wire main_rtio_core_outputs_selected163;
wire main_rtio_core_outputs_selected164;
wire main_rtio_core_outputs_selected165;
wire main_rtio_core_outputs_selected166;
wire main_rtio_core_outputs_selected167;
wire main_rtio_core_outputs_selected168;
wire main_rtio_core_outputs_selected169;
wire main_rtio_core_outputs_selected170;
wire main_rtio_core_outputs_selected171;
wire main_rtio_core_outputs_selected172;
wire main_rtio_core_outputs_selected173;
wire main_rtio_core_outputs_selected174;
wire main_rtio_core_outputs_selected175;
wire main_rtio_core_outputs_selected176;
wire main_rtio_core_outputs_selected177;
wire main_rtio_core_outputs_selected178;
wire main_rtio_core_outputs_selected179;
wire main_rtio_core_outputs_selected180;
wire main_rtio_core_outputs_selected181;
wire main_rtio_core_outputs_selected182;
wire main_rtio_core_outputs_selected183;
wire main_rtio_core_outputs_selected184;
wire main_rtio_core_outputs_selected185;
wire main_rtio_core_outputs_selected186;
wire main_rtio_core_outputs_selected187;
wire main_rtio_core_outputs_selected188;
wire main_rtio_core_outputs_selected189;
wire main_rtio_core_outputs_selected190;
wire main_rtio_core_outputs_selected191;
wire main_rtio_core_outputs_selected192;
wire main_rtio_core_outputs_selected193;
wire main_rtio_core_outputs_selected194;
wire main_rtio_core_outputs_selected195;
wire main_rtio_core_outputs_selected196;
wire main_rtio_core_outputs_selected197;
wire main_rtio_core_outputs_selected198;
wire main_rtio_core_outputs_selected199;
wire main_rtio_core_outputs_selected200;
wire main_rtio_core_outputs_selected201;
wire main_rtio_core_outputs_selected202;
wire main_rtio_core_outputs_selected203;
wire main_rtio_core_outputs_selected204;
wire main_rtio_core_outputs_selected205;
wire main_rtio_core_outputs_selected206;
wire main_rtio_core_outputs_selected207;
wire main_rtio_core_outputs_selected208;
wire main_rtio_core_outputs_selected209;
wire main_rtio_core_outputs_selected210;
wire main_rtio_core_outputs_selected211;
wire main_rtio_core_outputs_selected212;
wire main_rtio_core_outputs_selected213;
wire main_rtio_core_outputs_selected214;
wire main_rtio_core_outputs_selected215;
wire main_rtio_core_outputs_selected216;
wire main_rtio_core_outputs_selected217;
wire main_rtio_core_outputs_selected218;
wire main_rtio_core_outputs_selected219;
wire main_rtio_core_outputs_selected220;
wire main_rtio_core_outputs_selected221;
wire main_rtio_core_outputs_selected222;
wire main_rtio_core_outputs_selected223;
wire main_rtio_core_outputs_selected224;
wire main_rtio_core_outputs_selected225;
wire main_rtio_core_outputs_selected226;
wire main_rtio_core_outputs_selected227;
wire main_rtio_core_outputs_selected228;
wire main_rtio_core_outputs_selected229;
wire main_rtio_core_outputs_selected230;
wire main_rtio_core_outputs_selected231;
wire main_rtio_core_outputs_selected232;
wire main_rtio_core_outputs_selected233;
wire main_rtio_core_outputs_selected234;
wire main_rtio_core_outputs_selected235;
wire main_rtio_core_outputs_selected236;
wire main_rtio_core_outputs_selected237;
wire main_rtio_core_outputs_selected238;
wire main_rtio_core_outputs_selected239;
wire main_rtio_core_outputs_selected240;
wire main_rtio_core_outputs_selected241;
wire main_rtio_core_outputs_selected242;
wire main_rtio_core_outputs_selected243;
wire main_rtio_core_outputs_selected244;
wire main_rtio_core_outputs_selected245;
wire main_rtio_core_outputs_selected246;
wire main_rtio_core_outputs_selected247;
wire main_rtio_core_outputs_selected248;
wire main_rtio_core_outputs_selected249;
wire main_rtio_core_outputs_selected250;
wire main_rtio_core_outputs_selected251;
wire main_rtio_core_outputs_selected252;
wire main_rtio_core_outputs_selected253;
wire main_rtio_core_outputs_selected254;
wire main_rtio_core_outputs_selected255;
wire main_rtio_core_outputs_selected256;
wire main_rtio_core_outputs_selected257;
wire main_rtio_core_outputs_selected258;
wire main_rtio_core_outputs_selected259;
wire main_rtio_core_outputs_selected260;
wire main_rtio_core_outputs_selected261;
wire main_rtio_core_outputs_selected262;
wire main_rtio_core_outputs_selected263;
wire main_rtio_core_outputs_selected264;
wire main_rtio_core_outputs_selected265;
wire main_rtio_core_outputs_selected266;
wire main_rtio_core_outputs_selected267;
wire main_rtio_core_outputs_selected268;
wire main_rtio_core_outputs_selected269;
wire main_rtio_core_outputs_selected270;
wire main_rtio_core_outputs_selected271;
wire main_rtio_core_outputs_selected272;
wire main_rtio_core_outputs_selected273;
wire main_rtio_core_outputs_selected274;
wire main_rtio_core_outputs_selected275;
wire main_rtio_core_outputs_selected276;
wire main_rtio_core_outputs_selected277;
wire main_rtio_core_outputs_selected278;
wire main_rtio_core_outputs_selected279;
wire main_rtio_core_outputs_selected280;
wire main_rtio_core_outputs_selected281;
wire main_rtio_core_outputs_selected282;
wire main_rtio_core_outputs_selected283;
wire main_rtio_core_outputs_selected284;
wire main_rtio_core_outputs_selected285;
wire main_rtio_core_outputs_selected286;
wire main_rtio_core_outputs_selected287;
wire main_rtio_core_outputs_selected288;
wire main_rtio_core_outputs_selected289;
wire main_rtio_core_outputs_selected290;
wire main_rtio_core_outputs_selected291;
wire main_rtio_core_outputs_selected292;
wire main_rtio_core_outputs_selected293;
wire main_rtio_core_outputs_selected294;
wire main_rtio_core_outputs_selected295;
reg main_rtio_core_outputs_stb_r0 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r0 = 6'd0;
reg main_rtio_core_outputs_stb_r1 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r1 = 6'd0;
reg main_rtio_core_outputs_stb_r2 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r2 = 6'd0;
reg main_rtio_core_outputs_stb_r3 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r3 = 6'd0;
reg main_rtio_core_outputs_stb_r4 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r4 = 6'd0;
reg main_rtio_core_outputs_stb_r5 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r5 = 6'd0;
reg main_rtio_core_outputs_stb_r6 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r6 = 6'd0;
reg main_rtio_core_outputs_stb_r7 = 1'd0;
reg [5:0] main_rtio_core_outputs_channel_r7 = 6'd0;
reg main_rtio_core_inputs_i_ack = 1'd0;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_we;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_re;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
wire [64:0] main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
wire main_rtio_core_inputs_asyncfifo0_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
wire main_rtio_core_inputs_asyncfifo0_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo0_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo0_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo0_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo0_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo0_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo0_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo0_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo0_rdport_dat_r;
wire main_rtio_core_inputs_record0_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record0_fifo_in_timestamp;
wire main_rtio_core_inputs_record0_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record0_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io0;
wire main_rtio_core_inputs_blindtransfer0_i;
wire main_rtio_core_inputs_blindtransfer0_o;
wire main_rtio_core_inputs_blindtransfer0_ps_i;
wire main_rtio_core_inputs_blindtransfer0_ps_o;
reg main_rtio_core_inputs_blindtransfer0_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer0_blind = 1'd0;
wire main_rtio_core_inputs_selected0;
reg main_rtio_core_inputs_overflow0 = 1'd0;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_we;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_re;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
wire [64:0] main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
wire main_rtio_core_inputs_asyncfifo1_graycounter2_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
wire main_rtio_core_inputs_asyncfifo1_graycounter3_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo1_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo1_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo1_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo1_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo1_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo1_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo1_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo1_rdport_dat_r;
wire main_rtio_core_inputs_record1_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record1_fifo_in_timestamp;
wire main_rtio_core_inputs_record1_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record1_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io1;
wire main_rtio_core_inputs_blindtransfer1_i;
wire main_rtio_core_inputs_blindtransfer1_o;
wire main_rtio_core_inputs_blindtransfer1_ps_i;
wire main_rtio_core_inputs_blindtransfer1_ps_o;
reg main_rtio_core_inputs_blindtransfer1_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer1_blind = 1'd0;
wire main_rtio_core_inputs_selected1;
reg main_rtio_core_inputs_overflow1 = 1'd0;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_we;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_re;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
wire [64:0] main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
wire main_rtio_core_inputs_asyncfifo2_graycounter4_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
wire main_rtio_core_inputs_asyncfifo2_graycounter5_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo2_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo2_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo2_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo2_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo2_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo2_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo2_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo2_rdport_dat_r;
wire main_rtio_core_inputs_record2_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record2_fifo_in_timestamp;
wire main_rtio_core_inputs_record2_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record2_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io2;
wire main_rtio_core_inputs_blindtransfer2_i;
wire main_rtio_core_inputs_blindtransfer2_o;
wire main_rtio_core_inputs_blindtransfer2_ps_i;
wire main_rtio_core_inputs_blindtransfer2_ps_o;
reg main_rtio_core_inputs_blindtransfer2_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer2_blind = 1'd0;
wire main_rtio_core_inputs_selected2;
reg main_rtio_core_inputs_overflow2 = 1'd0;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_we;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_re;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
wire [64:0] main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
wire main_rtio_core_inputs_asyncfifo3_graycounter6_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
wire main_rtio_core_inputs_asyncfifo3_graycounter7_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo3_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo3_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo3_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo3_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo3_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo3_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo3_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo3_rdport_dat_r;
wire main_rtio_core_inputs_record3_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record3_fifo_in_timestamp;
wire main_rtio_core_inputs_record3_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record3_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io3;
wire main_rtio_core_inputs_blindtransfer3_i;
wire main_rtio_core_inputs_blindtransfer3_o;
wire main_rtio_core_inputs_blindtransfer3_ps_i;
wire main_rtio_core_inputs_blindtransfer3_ps_o;
reg main_rtio_core_inputs_blindtransfer3_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer3_blind = 1'd0;
wire main_rtio_core_inputs_selected3;
reg main_rtio_core_inputs_overflow3 = 1'd0;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_we;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_re;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
wire [64:0] main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
wire main_rtio_core_inputs_asyncfifo4_graycounter8_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
wire main_rtio_core_inputs_asyncfifo4_graycounter9_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo4_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo4_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo4_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo4_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo4_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo4_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo4_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo4_rdport_dat_r;
wire main_rtio_core_inputs_record4_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record4_fifo_in_timestamp;
wire main_rtio_core_inputs_record4_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record4_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io4;
wire main_rtio_core_inputs_blindtransfer4_i;
wire main_rtio_core_inputs_blindtransfer4_o;
wire main_rtio_core_inputs_blindtransfer4_ps_i;
wire main_rtio_core_inputs_blindtransfer4_ps_o;
reg main_rtio_core_inputs_blindtransfer4_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer4_blind = 1'd0;
wire main_rtio_core_inputs_selected4;
reg main_rtio_core_inputs_overflow4 = 1'd0;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_we;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_re;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
wire [64:0] main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
wire main_rtio_core_inputs_asyncfifo5_graycounter10_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
wire main_rtio_core_inputs_asyncfifo5_graycounter11_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo5_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo5_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo5_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo5_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo5_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo5_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo5_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo5_rdport_dat_r;
wire main_rtio_core_inputs_record5_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record5_fifo_in_timestamp;
wire main_rtio_core_inputs_record5_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record5_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io5;
wire main_rtio_core_inputs_blindtransfer5_i;
wire main_rtio_core_inputs_blindtransfer5_o;
wire main_rtio_core_inputs_blindtransfer5_ps_i;
wire main_rtio_core_inputs_blindtransfer5_ps_o;
reg main_rtio_core_inputs_blindtransfer5_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer5_blind = 1'd0;
wire main_rtio_core_inputs_selected5;
reg main_rtio_core_inputs_overflow5 = 1'd0;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_we;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_re;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
wire [64:0] main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
wire main_rtio_core_inputs_asyncfifo6_graycounter12_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
wire main_rtio_core_inputs_asyncfifo6_graycounter13_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo6_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo6_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo6_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo6_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo6_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo6_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo6_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo6_rdport_dat_r;
wire main_rtio_core_inputs_record6_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record6_fifo_in_timestamp;
wire main_rtio_core_inputs_record6_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record6_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io6;
wire main_rtio_core_inputs_blindtransfer6_i;
wire main_rtio_core_inputs_blindtransfer6_o;
wire main_rtio_core_inputs_blindtransfer6_ps_i;
wire main_rtio_core_inputs_blindtransfer6_ps_o;
reg main_rtio_core_inputs_blindtransfer6_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer6_blind = 1'd0;
wire main_rtio_core_inputs_selected6;
reg main_rtio_core_inputs_overflow6 = 1'd0;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_we;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_re;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo7_asyncfifo7_din;
wire [64:0] main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout;
wire main_rtio_core_inputs_asyncfifo7_graycounter14_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary;
wire main_rtio_core_inputs_asyncfifo7_graycounter15_ce;
(* dont_touch = "true" *) reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q = 7'd0;
wire [6:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_next;
reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary = 7'd0;
reg [6:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary;
wire [6:0] main_rtio_core_inputs_asyncfifo7_produce_rdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo7_consume_wdomain;
wire [5:0] main_rtio_core_inputs_asyncfifo7_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo7_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo7_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo7_wrport_dat_w;
wire [5:0] main_rtio_core_inputs_asyncfifo7_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo7_rdport_dat_r;
wire main_rtio_core_inputs_record7_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record7_fifo_in_timestamp;
wire main_rtio_core_inputs_record7_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record7_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io7;
wire main_rtio_core_inputs_blindtransfer7_i;
wire main_rtio_core_inputs_blindtransfer7_o;
wire main_rtio_core_inputs_blindtransfer7_ps_i;
wire main_rtio_core_inputs_blindtransfer7_ps_o;
reg main_rtio_core_inputs_blindtransfer7_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer7_blind = 1'd0;
wire main_rtio_core_inputs_selected7;
reg main_rtio_core_inputs_overflow7 = 1'd0;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_we;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_re;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo8_asyncfifo8_din;
wire [31:0] main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout;
wire main_rtio_core_inputs_asyncfifo8_graycounter16_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary;
wire main_rtio_core_inputs_asyncfifo8_graycounter17_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary;
wire [2:0] main_rtio_core_inputs_asyncfifo8_produce_rdomain;
wire [2:0] main_rtio_core_inputs_asyncfifo8_consume_wdomain;
wire [1:0] main_rtio_core_inputs_asyncfifo8_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo8_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo8_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo8_wrport_dat_w;
wire [1:0] main_rtio_core_inputs_asyncfifo8_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo8_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record8_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record8_fifo_out_data;
wire main_rtio_core_inputs_overflow_io8;
wire main_rtio_core_inputs_blindtransfer8_i;
wire main_rtio_core_inputs_blindtransfer8_o;
wire main_rtio_core_inputs_blindtransfer8_ps_i;
wire main_rtio_core_inputs_blindtransfer8_ps_o;
reg main_rtio_core_inputs_blindtransfer8_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer8_blind = 1'd0;
wire main_rtio_core_inputs_selected8;
reg main_rtio_core_inputs_overflow8 = 1'd0;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_we;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_re;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo9_asyncfifo9_din;
wire [31:0] main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout;
wire main_rtio_core_inputs_asyncfifo9_graycounter18_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary;
wire main_rtio_core_inputs_asyncfifo9_graycounter19_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary;
wire [2:0] main_rtio_core_inputs_asyncfifo9_produce_rdomain;
wire [2:0] main_rtio_core_inputs_asyncfifo9_consume_wdomain;
wire [1:0] main_rtio_core_inputs_asyncfifo9_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo9_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo9_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo9_wrport_dat_w;
wire [1:0] main_rtio_core_inputs_asyncfifo9_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo9_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record9_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record9_fifo_out_data;
wire main_rtio_core_inputs_overflow_io9;
wire main_rtio_core_inputs_blindtransfer9_i;
wire main_rtio_core_inputs_blindtransfer9_o;
wire main_rtio_core_inputs_blindtransfer9_ps_i;
wire main_rtio_core_inputs_blindtransfer9_ps_o;
reg main_rtio_core_inputs_blindtransfer9_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer9_blind = 1'd0;
wire main_rtio_core_inputs_selected9;
reg main_rtio_core_inputs_overflow9 = 1'd0;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_we;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_re;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo10_asyncfifo10_din;
wire [31:0] main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout;
wire main_rtio_core_inputs_asyncfifo10_graycounter20_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary;
wire main_rtio_core_inputs_asyncfifo10_graycounter21_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary;
wire [2:0] main_rtio_core_inputs_asyncfifo10_produce_rdomain;
wire [2:0] main_rtio_core_inputs_asyncfifo10_consume_wdomain;
wire [1:0] main_rtio_core_inputs_asyncfifo10_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo10_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo10_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo10_wrport_dat_w;
wire [1:0] main_rtio_core_inputs_asyncfifo10_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo10_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record10_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record10_fifo_out_data;
wire main_rtio_core_inputs_overflow_io10;
wire main_rtio_core_inputs_blindtransfer10_i;
wire main_rtio_core_inputs_blindtransfer10_o;
wire main_rtio_core_inputs_blindtransfer10_ps_i;
wire main_rtio_core_inputs_blindtransfer10_ps_o;
reg main_rtio_core_inputs_blindtransfer10_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer10_blind = 1'd0;
wire main_rtio_core_inputs_selected10;
reg main_rtio_core_inputs_overflow10 = 1'd0;
wire [1:0] main_rtio_core_inputs_i_status_raw;
reg [63:0] main_rtio_core_inputs_input_timeout = 64'd0;
reg main_rtio_core_inputs_input_pending = 1'd0;
wire main_rtio_core_o_collision_sync_i;
wire main_rtio_core_o_collision_sync_o;
wire [15:0] main_rtio_core_o_collision_sync_data_i;
wire [15:0] main_rtio_core_o_collision_sync_data_o;
wire main_rtio_core_o_collision_sync_ps_i;
wire main_rtio_core_o_collision_sync_ps_o;
reg main_rtio_core_o_collision_sync_ps_toggle_i = 1'd0;
wire main_rtio_core_o_collision_sync_ps_toggle_o;
reg main_rtio_core_o_collision_sync_ps_toggle_o_r = 1'd0;
wire main_rtio_core_o_collision_sync_ps_ack_i;
wire main_rtio_core_o_collision_sync_ps_ack_o;
reg main_rtio_core_o_collision_sync_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_o_collision_sync_ps_ack_toggle_o;
reg main_rtio_core_o_collision_sync_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_o_collision_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_rtio_core_o_collision_sync_bxfer_data = 16'd0;
wire main_rtio_core_o_busy_sync_i;
wire main_rtio_core_o_busy_sync_o;
wire [15:0] main_rtio_core_o_busy_sync_data_i;
wire [15:0] main_rtio_core_o_busy_sync_data_o;
wire main_rtio_core_o_busy_sync_ps_i;
wire main_rtio_core_o_busy_sync_ps_o;
reg main_rtio_core_o_busy_sync_ps_toggle_i = 1'd0;
wire main_rtio_core_o_busy_sync_ps_toggle_o;
reg main_rtio_core_o_busy_sync_ps_toggle_o_r = 1'd0;
wire main_rtio_core_o_busy_sync_ps_ack_i;
wire main_rtio_core_o_busy_sync_ps_ack_o;
reg main_rtio_core_o_busy_sync_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_o_busy_sync_ps_ack_toggle_o;
reg main_rtio_core_o_busy_sync_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_o_busy_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_rtio_core_o_busy_sync_bxfer_data = 16'd0;
reg main_rtio_core_o_collision = 1'd0;
reg main_rtio_core_o_busy = 1'd0;
reg main_rtio_core_o_sequence_error = 1'd0;
reg [31:0] main_rtio_target_storage_full = 32'd0;
wire [31:0] main_rtio_target_storage;
reg main_rtio_target_re = 1'd0;
wire main_rtio_now_hi_re;
wire [31:0] main_rtio_now_hi_r;
wire [31:0] main_rtio_now_hi_w;
wire main_rtio_now_lo_re;
wire [31:0] main_rtio_now_lo_r;
wire [31:0] main_rtio_now_lo_w;
reg [511:0] main_rtio_o_data_storage_full = 512'd0;
wire [511:0] main_rtio_o_data_storage;
reg main_rtio_o_data_re = 1'd0;
wire main_rtio_o_data_we;
wire [511:0] main_rtio_o_data_dat_w;
wire [2:0] main_rtio_o_status_status;
reg [63:0] main_rtio_i_timeout_storage_full = 64'd0;
wire [63:0] main_rtio_i_timeout_storage;
reg main_rtio_i_timeout_re = 1'd0;
wire [31:0] main_rtio_i_data_status;
wire [63:0] main_rtio_i_timestamp_status;
wire [3:0] main_rtio_i_status_status;
wire main_rtio_i_overflow_reset_re;
wire main_rtio_i_overflow_reset_r;
reg main_rtio_i_overflow_reset_w = 1'd0;
reg [63:0] main_rtio_counter_status = 64'd0;
wire main_rtio_counter_update_re;
wire main_rtio_counter_update_r;
reg main_rtio_counter_update_w = 1'd0;
reg [1:0] main_rtio_cri_cmd;
wire [23:0] main_rtio_cri_chan_sel;
wire [63:0] main_rtio_cri_o_timestamp;
wire [511:0] main_rtio_cri_o_data;
wire [7:0] main_rtio_cri_o_address;
wire [2:0] main_rtio_cri_o_status;
wire main_rtio_cri_o_buffer_space_valid;
wire [15:0] main_rtio_cri_o_buffer_space;
wire [63:0] main_rtio_cri_i_timeout;
wire [31:0] main_rtio_cri_i_data;
wire [63:0] main_rtio_cri_i_timestamp;
wire [3:0] main_rtio_cri_i_status;
reg [31:0] main_rtio_now_hi_backing = 32'd0;
reg [63:0] main_rtio_now = 64'd0;
wire [29:0] main_genericstandalone_interface0_bus_adr;
reg [127:0] main_genericstandalone_interface0_bus_dat_w = 128'd0;
wire [127:0] main_genericstandalone_interface0_bus_dat_r;
reg [15:0] main_genericstandalone_interface0_bus_sel = 16'd0;
wire main_genericstandalone_interface0_bus_cyc;
wire main_genericstandalone_interface0_bus_stb;
wire main_genericstandalone_interface0_bus_ack;
reg main_genericstandalone_interface0_bus_we = 1'd0;
reg [2:0] main_genericstandalone_interface0_bus_cti = 3'd0;
reg [1:0] main_genericstandalone_interface0_bus_bte = 2'd0;
wire main_genericstandalone_interface0_bus_err;
wire main_dma_enable_enable_re;
wire main_dma_enable_enable_r;
reg main_dma_enable_enable_w;
reg main_dma_flow_enable;
reg main_dma_dma_sink_stb = 1'd0;
wire main_dma_dma_sink_ack;
reg main_dma_dma_sink_eop = 1'd0;
reg [29:0] main_dma_dma_sink_payload_address = 30'd0;
wire main_dma_dma_source_stb;
wire main_dma_dma_source_ack;
reg main_dma_dma_source_eop = 1'd0;
reg [127:0] main_dma_dma_source_payload_data = 128'd0;
wire main_dma_dma_bus_stb;
reg main_dma_dma_data_reg_loaded = 1'd0;
reg [33:0] main_dma_dma_storage_full = 34'd0;
wire [29:0] main_dma_dma_storage;
reg main_dma_dma_re = 1'd0;
reg main_dma_dma_enable_r = 1'd0;
wire main_dma_rawslicer_sink_stb;
reg main_dma_rawslicer_sink_ack;
wire main_dma_rawslicer_sink_eop;
wire [127:0] main_dma_rawslicer_sink_payload_data;
wire [615:0] main_dma_rawslicer_source;
reg main_dma_rawslicer_source_stb;
reg [6:0] main_dma_rawslicer_source_consume;
reg main_dma_rawslicer_flush;
reg main_dma_rawslicer_flush_done;
reg [735:0] main_dma_rawslicer_buf = 736'd0;
reg [6:0] main_dma_rawslicer_level = 7'd0;
reg [6:0] main_dma_rawslicer_next_level;
reg main_dma_rawslicer_load_buf;
reg main_dma_rawslicer_shift_buf;
reg main_dma_reset = 1'd0;
reg main_dma_record_converter_source_stb;
wire main_dma_record_converter_source_ack;
reg main_dma_record_converter_source_eop;
reg [7:0] main_dma_record_converter_source_payload_length = 8'd0;
wire [23:0] main_dma_record_converter_source_payload_channel;
wire [63:0] main_dma_record_converter_source_payload_timestamp;
wire [7:0] main_dma_record_converter_source_payload_address;
reg [511:0] main_dma_record_converter_source_payload_data;
reg main_dma_record_converter_end_marker_found;
reg main_dma_record_converter_flush;
wire [7:0] main_dma_record_converter_record_raw_length;
wire [23:0] main_dma_record_converter_record_raw_channel;
wire [63:0] main_dma_record_converter_record_raw_timestamp;
wire [7:0] main_dma_record_converter_record_raw_address;
wire [511:0] main_dma_record_converter_record_raw_data;
reg [63:0] main_dma_time_offset_storage_full = 64'd0;
wire [63:0] main_dma_time_offset_storage;
reg main_dma_time_offset_re = 1'd0;
reg main_dma_time_offset_source_stb = 1'd0;
wire main_dma_time_offset_source_ack;
reg main_dma_time_offset_source_eop = 1'd0;
reg [7:0] main_dma_time_offset_source_payload_length = 8'd0;
reg [23:0] main_dma_time_offset_source_payload_channel = 24'd0;
reg [63:0] main_dma_time_offset_source_payload_timestamp = 64'd0;
reg [7:0] main_dma_time_offset_source_payload_address = 8'd0;
reg [511:0] main_dma_time_offset_source_payload_data = 512'd0;
wire main_dma_time_offset_sink_stb;
wire main_dma_time_offset_sink_ack;
wire main_dma_time_offset_sink_eop;
wire [7:0] main_dma_time_offset_sink_payload_length;
wire [23:0] main_dma_time_offset_sink_payload_channel;
wire [63:0] main_dma_time_offset_sink_payload_timestamp;
wire [7:0] main_dma_time_offset_sink_payload_address;
wire [511:0] main_dma_time_offset_sink_payload_data;
wire main_dma_cri_master_error_re;
wire [1:0] main_dma_cri_master_error_r;
reg [1:0] main_dma_cri_master_error_w = 2'd0;
reg [23:0] main_dma_cri_master_error_channel_status = 24'd0;
reg [63:0] main_dma_cri_master_error_timestamp_status = 64'd0;
reg [15:0] main_dma_cri_master_error_address_status = 16'd0;
wire main_dma_cri_master_sink_stb;
reg main_dma_cri_master_sink_ack;
wire main_dma_cri_master_sink_eop;
wire [7:0] main_dma_cri_master_sink_payload_length;
wire [23:0] main_dma_cri_master_sink_payload_channel;
wire [63:0] main_dma_cri_master_sink_payload_timestamp;
wire [7:0] main_dma_cri_master_sink_payload_address;
wire [511:0] main_dma_cri_master_sink_payload_data;
reg [1:0] main_dma_cri_master_cri_cmd;
wire [23:0] main_dma_cri_master_cri_chan_sel;
wire [63:0] main_dma_cri_master_cri_o_timestamp;
wire [511:0] main_dma_cri_master_cri_o_data;
wire [7:0] main_dma_cri_master_cri_o_address;
wire [2:0] main_dma_cri_master_cri_o_status;
wire main_dma_cri_master_cri_o_buffer_space_valid;
wire [15:0] main_dma_cri_master_cri_o_buffer_space;
reg [63:0] main_dma_cri_master_cri_i_timeout = 64'd0;
wire [31:0] main_dma_cri_master_cri_i_data;
wire [63:0] main_dma_cri_master_cri_i_timestamp;
wire [3:0] main_dma_cri_master_cri_i_status;
reg main_dma_cri_master_busy;
reg main_dma_cri_master_underflow_trigger;
reg main_dma_cri_master_link_error_trigger;
wire [29:0] main_genericstandalone_csrbank0_bus_adr;
wire [31:0] main_genericstandalone_csrbank0_bus_dat_w;
reg [31:0] main_genericstandalone_csrbank0_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_csrbank0_bus_sel;
wire main_genericstandalone_csrbank0_bus_cyc;
wire main_genericstandalone_csrbank0_bus_stb;
reg main_genericstandalone_csrbank0_bus_ack = 1'd0;
wire main_genericstandalone_csrbank0_bus_we;
wire [2:0] main_genericstandalone_csrbank0_bus_cti;
wire [1:0] main_genericstandalone_csrbank0_bus_bte;
reg main_genericstandalone_csrbank0_bus_err = 1'd0;
wire main_genericstandalone_csrbank0_target0_re;
wire [31:0] main_genericstandalone_csrbank0_target0_r;
wire [31:0] main_genericstandalone_csrbank0_target0_w;
wire main_genericstandalone_csrbank0_o_data15_re;
wire [31:0] main_genericstandalone_csrbank0_o_data15_r;
wire [31:0] main_genericstandalone_csrbank0_o_data15_w;
wire main_genericstandalone_csrbank0_o_data14_re;
wire [31:0] main_genericstandalone_csrbank0_o_data14_r;
wire [31:0] main_genericstandalone_csrbank0_o_data14_w;
wire main_genericstandalone_csrbank0_o_data13_re;
wire [31:0] main_genericstandalone_csrbank0_o_data13_r;
wire [31:0] main_genericstandalone_csrbank0_o_data13_w;
wire main_genericstandalone_csrbank0_o_data12_re;
wire [31:0] main_genericstandalone_csrbank0_o_data12_r;
wire [31:0] main_genericstandalone_csrbank0_o_data12_w;
wire main_genericstandalone_csrbank0_o_data11_re;
wire [31:0] main_genericstandalone_csrbank0_o_data11_r;
wire [31:0] main_genericstandalone_csrbank0_o_data11_w;
wire main_genericstandalone_csrbank0_o_data10_re;
wire [31:0] main_genericstandalone_csrbank0_o_data10_r;
wire [31:0] main_genericstandalone_csrbank0_o_data10_w;
wire main_genericstandalone_csrbank0_o_data9_re;
wire [31:0] main_genericstandalone_csrbank0_o_data9_r;
wire [31:0] main_genericstandalone_csrbank0_o_data9_w;
wire main_genericstandalone_csrbank0_o_data8_re;
wire [31:0] main_genericstandalone_csrbank0_o_data8_r;
wire [31:0] main_genericstandalone_csrbank0_o_data8_w;
wire main_genericstandalone_csrbank0_o_data7_re;
wire [31:0] main_genericstandalone_csrbank0_o_data7_r;
wire [31:0] main_genericstandalone_csrbank0_o_data7_w;
wire main_genericstandalone_csrbank0_o_data6_re;
wire [31:0] main_genericstandalone_csrbank0_o_data6_r;
wire [31:0] main_genericstandalone_csrbank0_o_data6_w;
wire main_genericstandalone_csrbank0_o_data5_re;
wire [31:0] main_genericstandalone_csrbank0_o_data5_r;
wire [31:0] main_genericstandalone_csrbank0_o_data5_w;
wire main_genericstandalone_csrbank0_o_data4_re;
wire [31:0] main_genericstandalone_csrbank0_o_data4_r;
wire [31:0] main_genericstandalone_csrbank0_o_data4_w;
wire main_genericstandalone_csrbank0_o_data3_re;
wire [31:0] main_genericstandalone_csrbank0_o_data3_r;
wire [31:0] main_genericstandalone_csrbank0_o_data3_w;
wire main_genericstandalone_csrbank0_o_data2_re;
wire [31:0] main_genericstandalone_csrbank0_o_data2_r;
wire [31:0] main_genericstandalone_csrbank0_o_data2_w;
wire main_genericstandalone_csrbank0_o_data1_re;
wire [31:0] main_genericstandalone_csrbank0_o_data1_r;
wire [31:0] main_genericstandalone_csrbank0_o_data1_w;
wire main_genericstandalone_csrbank0_o_data0_re;
wire [31:0] main_genericstandalone_csrbank0_o_data0_r;
wire [31:0] main_genericstandalone_csrbank0_o_data0_w;
wire main_genericstandalone_csrbank0_o_status_re;
wire [2:0] main_genericstandalone_csrbank0_o_status_r;
wire [2:0] main_genericstandalone_csrbank0_o_status_w;
wire main_genericstandalone_csrbank0_i_timeout1_re;
wire [31:0] main_genericstandalone_csrbank0_i_timeout1_r;
wire [31:0] main_genericstandalone_csrbank0_i_timeout1_w;
wire main_genericstandalone_csrbank0_i_timeout0_re;
wire [31:0] main_genericstandalone_csrbank0_i_timeout0_r;
wire [31:0] main_genericstandalone_csrbank0_i_timeout0_w;
wire main_genericstandalone_csrbank0_i_data_re;
wire [31:0] main_genericstandalone_csrbank0_i_data_r;
wire [31:0] main_genericstandalone_csrbank0_i_data_w;
wire main_genericstandalone_csrbank0_i_timestamp1_re;
wire [31:0] main_genericstandalone_csrbank0_i_timestamp1_r;
wire [31:0] main_genericstandalone_csrbank0_i_timestamp1_w;
wire main_genericstandalone_csrbank0_i_timestamp0_re;
wire [31:0] main_genericstandalone_csrbank0_i_timestamp0_r;
wire [31:0] main_genericstandalone_csrbank0_i_timestamp0_w;
wire main_genericstandalone_csrbank0_i_status_re;
wire [3:0] main_genericstandalone_csrbank0_i_status_r;
wire [3:0] main_genericstandalone_csrbank0_i_status_w;
wire main_genericstandalone_csrbank0_counter1_re;
wire [31:0] main_genericstandalone_csrbank0_counter1_r;
wire [31:0] main_genericstandalone_csrbank0_counter1_w;
wire main_genericstandalone_csrbank0_counter0_re;
wire [31:0] main_genericstandalone_csrbank0_counter0_r;
wire [31:0] main_genericstandalone_csrbank0_counter0_w;
wire [29:0] main_genericstandalone_csrbank1_bus_adr;
wire [31:0] main_genericstandalone_csrbank1_bus_dat_w;
reg [31:0] main_genericstandalone_csrbank1_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_csrbank1_bus_sel;
wire main_genericstandalone_csrbank1_bus_cyc;
wire main_genericstandalone_csrbank1_bus_stb;
reg main_genericstandalone_csrbank1_bus_ack = 1'd0;
wire main_genericstandalone_csrbank1_bus_we;
wire [2:0] main_genericstandalone_csrbank1_bus_cti;
wire [1:0] main_genericstandalone_csrbank1_bus_bte;
reg main_genericstandalone_csrbank1_bus_err = 1'd0;
wire main_genericstandalone_csrbank1_base_address1_re;
wire [1:0] main_genericstandalone_csrbank1_base_address1_r;
wire [1:0] main_genericstandalone_csrbank1_base_address1_w;
wire main_genericstandalone_csrbank1_base_address0_re;
wire [31:0] main_genericstandalone_csrbank1_base_address0_r;
wire [31:0] main_genericstandalone_csrbank1_base_address0_w;
wire main_genericstandalone_csrbank1_time_offset1_re;
wire [31:0] main_genericstandalone_csrbank1_time_offset1_r;
wire [31:0] main_genericstandalone_csrbank1_time_offset1_w;
wire main_genericstandalone_csrbank1_time_offset0_re;
wire [31:0] main_genericstandalone_csrbank1_time_offset0_r;
wire [31:0] main_genericstandalone_csrbank1_time_offset0_w;
wire main_genericstandalone_csrbank1_error_channel_re;
wire [23:0] main_genericstandalone_csrbank1_error_channel_r;
wire [23:0] main_genericstandalone_csrbank1_error_channel_w;
wire main_genericstandalone_csrbank1_error_timestamp1_re;
wire [31:0] main_genericstandalone_csrbank1_error_timestamp1_r;
wire [31:0] main_genericstandalone_csrbank1_error_timestamp1_w;
wire main_genericstandalone_csrbank1_error_timestamp0_re;
wire [31:0] main_genericstandalone_csrbank1_error_timestamp0_r;
wire [31:0] main_genericstandalone_csrbank1_error_timestamp0_w;
wire main_genericstandalone_csrbank1_error_address_re;
wire [15:0] main_genericstandalone_csrbank1_error_address_r;
wire [15:0] main_genericstandalone_csrbank1_error_address_w;
wire [1:0] main_cri_con_shared_cmd;
wire [23:0] main_cri_con_shared_chan_sel;
wire [63:0] main_cri_con_shared_o_timestamp;
wire [511:0] main_cri_con_shared_o_data;
wire [7:0] main_cri_con_shared_o_address;
reg [2:0] main_cri_con_shared_o_status;
reg main_cri_con_shared_o_buffer_space_valid;
reg [15:0] main_cri_con_shared_o_buffer_space;
wire [63:0] main_cri_con_shared_i_timeout;
reg [31:0] main_cri_con_shared_i_data;
reg [63:0] main_cri_con_shared_i_timestamp;
reg [3:0] main_cri_con_shared_i_status;
reg [1:0] main_cri_con_storage_full = 2'd0;
wire [1:0] main_cri_con_storage;
reg main_cri_con_re = 1'd0;
reg main_cri_con_selected = 1'd0;
wire [29:0] main_genericstandalone_csrbank2_bus_adr;
wire [31:0] main_genericstandalone_csrbank2_bus_dat_w;
reg [31:0] main_genericstandalone_csrbank2_bus_dat_r = 32'd0;
wire [3:0] main_genericstandalone_csrbank2_bus_sel;
wire main_genericstandalone_csrbank2_bus_cyc;
wire main_genericstandalone_csrbank2_bus_stb;
reg main_genericstandalone_csrbank2_bus_ack = 1'd0;
wire main_genericstandalone_csrbank2_bus_we;
wire [2:0] main_genericstandalone_csrbank2_bus_cti;
wire [1:0] main_genericstandalone_csrbank2_bus_bte;
reg main_genericstandalone_csrbank2_bus_err = 1'd0;
wire main_genericstandalone_csrbank2_selected0_re;
wire [1:0] main_genericstandalone_csrbank2_selected0_r;
wire [1:0] main_genericstandalone_csrbank2_selected0_w;
reg [5:0] main_mon_chan_sel_storage_full = 6'd0;
wire [5:0] main_mon_chan_sel_storage;
reg main_mon_chan_sel_re = 1'd0;
reg main_mon_probe_sel_storage_full = 1'd0;
wire main_mon_probe_sel_storage;
reg main_mon_probe_sel_re = 1'd0;
wire main_mon_value_update_re;
wire main_mon_value_update_r;
reg main_mon_value_update_w = 1'd0;
reg main_mon_status = 1'd0;
wire main_mon_bussynchronizer0_i;
wire main_mon_bussynchronizer0_o;
wire main_mon_bussynchronizer1_i;
wire main_mon_bussynchronizer1_o;
wire main_mon_bussynchronizer2_i;
wire main_mon_bussynchronizer2_o;
wire main_mon_bussynchronizer3_i;
wire main_mon_bussynchronizer3_o;
wire main_mon_bussynchronizer4_i;
wire main_mon_bussynchronizer4_o;
wire main_mon_bussynchronizer5_i;
wire main_mon_bussynchronizer5_o;
wire main_mon_bussynchronizer6_i;
wire main_mon_bussynchronizer6_o;
wire main_mon_bussynchronizer7_i;
wire main_mon_bussynchronizer7_o;
wire main_mon_bussynchronizer8_i;
wire main_mon_bussynchronizer8_o;
wire main_mon_bussynchronizer9_i;
wire main_mon_bussynchronizer9_o;
wire main_mon_bussynchronizer10_i;
wire main_mon_bussynchronizer10_o;
wire main_mon_bussynchronizer11_i;
wire main_mon_bussynchronizer11_o;
wire main_mon_bussynchronizer12_i;
wire main_mon_bussynchronizer12_o;
wire main_mon_bussynchronizer13_i;
wire main_mon_bussynchronizer13_o;
wire main_mon_bussynchronizer14_i;
wire main_mon_bussynchronizer14_o;
wire main_mon_bussynchronizer15_i;
wire main_mon_bussynchronizer15_o;
wire main_mon_bussynchronizer16_i;
wire main_mon_bussynchronizer16_o;
wire main_mon_bussynchronizer17_i;
wire main_mon_bussynchronizer17_o;
wire main_mon_bussynchronizer18_i;
wire main_mon_bussynchronizer18_o;
wire main_mon_bussynchronizer19_i;
wire main_mon_bussynchronizer19_o;
wire main_mon_bussynchronizer20_i;
wire main_mon_bussynchronizer20_o;
wire main_mon_bussynchronizer21_i;
wire main_mon_bussynchronizer21_o;
wire main_mon_bussynchronizer22_i;
wire main_mon_bussynchronizer22_o;
wire main_mon_bussynchronizer23_i;
wire main_mon_bussynchronizer23_o;
wire main_mon_bussynchronizer24_i;
wire main_mon_bussynchronizer24_o;
wire main_mon_bussynchronizer25_i;
wire main_mon_bussynchronizer25_o;
wire main_mon_bussynchronizer26_i;
wire main_mon_bussynchronizer26_o;
wire main_mon_bussynchronizer27_i;
wire main_mon_bussynchronizer27_o;
wire main_mon_bussynchronizer28_i;
wire main_mon_bussynchronizer28_o;
wire main_mon_bussynchronizer29_i;
wire main_mon_bussynchronizer29_o;
wire main_mon_bussynchronizer30_i;
wire main_mon_bussynchronizer30_o;
wire main_mon_bussynchronizer31_i;
wire main_mon_bussynchronizer31_o;
wire main_mon_bussynchronizer32_i;
wire main_mon_bussynchronizer32_o;
wire main_mon_bussynchronizer33_i;
wire main_mon_bussynchronizer33_o;
wire main_mon_bussynchronizer34_i;
wire main_mon_bussynchronizer34_o;
wire main_mon_bussynchronizer35_i;
wire main_mon_bussynchronizer35_o;
wire main_mon_bussynchronizer36_i;
wire main_mon_bussynchronizer36_o;
wire main_mon_bussynchronizer37_i;
wire main_mon_bussynchronizer37_o;
wire main_mon_bussynchronizer38_i;
wire main_mon_bussynchronizer38_o;
wire main_mon_bussynchronizer39_i;
wire main_mon_bussynchronizer39_o;
wire main_mon_bussynchronizer40_i;
wire main_mon_bussynchronizer40_o;
reg [5:0] main_inj_chan_sel_storage_full = 6'd0;
wire [5:0] main_inj_chan_sel_storage;
reg main_inj_chan_sel_re = 1'd0;
reg [1:0] main_inj_override_sel_storage_full = 2'd0;
wire [1:0] main_inj_override_sel_storage;
reg main_inj_override_sel_re = 1'd0;
wire main_inj_value_re;
wire main_inj_value_r;
wire main_inj_value_w;
reg main_inj_o_sys0 = 1'd0;
reg main_inj_o_sys1 = 1'd0;
reg main_inj_o_sys2 = 1'd0;
reg main_inj_o_sys3 = 1'd0;
reg main_inj_o_sys4 = 1'd0;
reg main_inj_o_sys5 = 1'd0;
reg main_inj_o_sys6 = 1'd0;
reg main_inj_o_sys7 = 1'd0;
reg main_inj_o_sys8 = 1'd0;
reg main_inj_o_sys9 = 1'd0;
reg main_inj_o_sys10 = 1'd0;
reg main_inj_o_sys11 = 1'd0;
reg main_inj_o_sys12 = 1'd0;
reg main_inj_o_sys13 = 1'd0;
reg main_inj_o_sys14 = 1'd0;
reg main_inj_o_sys15 = 1'd0;
reg main_inj_o_sys16 = 1'd0;
reg main_inj_o_sys17 = 1'd0;
reg main_inj_o_sys18 = 1'd0;
reg main_inj_o_sys19 = 1'd0;
reg main_inj_o_sys20 = 1'd0;
reg main_inj_o_sys21 = 1'd0;
reg main_inj_o_sys22 = 1'd0;
reg main_inj_o_sys23 = 1'd0;
reg main_inj_o_sys24 = 1'd0;
reg main_inj_o_sys25 = 1'd0;
reg main_inj_o_sys26 = 1'd0;
reg main_inj_o_sys27 = 1'd0;
reg main_inj_o_sys28 = 1'd0;
reg main_inj_o_sys29 = 1'd0;
reg main_inj_o_sys30 = 1'd0;
reg main_inj_o_sys31 = 1'd0;
reg main_inj_o_sys32 = 1'd0;
reg main_inj_o_sys33 = 1'd0;
reg main_inj_o_sys34 = 1'd0;
reg main_inj_o_sys35 = 1'd0;
reg main_inj_o_sys36 = 1'd0;
reg main_inj_o_sys37 = 1'd0;
reg main_inj_o_sys38 = 1'd0;
reg main_inj_o_sys39 = 1'd0;
reg main_inj_o_sys40 = 1'd0;
reg main_inj_o_sys41 = 1'd0;
reg main_inj_o_sys42 = 1'd0;
reg main_inj_o_sys43 = 1'd0;
reg main_inj_o_sys44 = 1'd0;
reg main_inj_o_sys45 = 1'd0;
reg main_inj_o_sys46 = 1'd0;
reg main_inj_o_sys47 = 1'd0;
reg main_inj_o_sys48 = 1'd0;
reg main_inj_o_sys49 = 1'd0;
reg main_inj_o_sys50 = 1'd0;
reg main_inj_o_sys51 = 1'd0;
reg main_inj_o_sys52 = 1'd0;
reg main_inj_o_sys53 = 1'd0;
reg main_inj_o_sys54 = 1'd0;
reg main_inj_o_sys55 = 1'd0;
reg main_inj_o_sys56 = 1'd0;
reg main_inj_o_sys57 = 1'd0;
reg main_inj_o_sys58 = 1'd0;
reg main_inj_o_sys59 = 1'd0;
reg main_inj_o_sys60 = 1'd0;
reg main_inj_o_sys61 = 1'd0;
reg main_inj_o_sys62 = 1'd0;
reg main_inj_o_sys63 = 1'd0;
reg main_inj_o_sys64 = 1'd0;
reg main_inj_o_sys65 = 1'd0;
reg main_inj_o_sys66 = 1'd0;
reg main_inj_o_sys67 = 1'd0;
reg main_inj_o_sys68 = 1'd0;
reg main_inj_o_sys69 = 1'd0;
reg main_inj_o_sys70 = 1'd0;
reg main_inj_o_sys71 = 1'd0;
reg main_inj_o_sys72 = 1'd0;
reg main_inj_o_sys73 = 1'd0;
reg [29:0] main_genericstandalone_interface1_bus_adr = 30'd0;
wire [127:0] main_genericstandalone_interface1_bus_dat_w;
wire [127:0] main_genericstandalone_interface1_bus_dat_r;
wire [15:0] main_genericstandalone_interface1_bus_sel;
wire main_genericstandalone_interface1_bus_cyc;
wire main_genericstandalone_interface1_bus_stb;
wire main_genericstandalone_interface1_bus_ack;
wire main_genericstandalone_interface1_bus_we;
reg [2:0] main_genericstandalone_interface1_bus_cti = 3'd0;
reg [1:0] main_genericstandalone_interface1_bus_bte = 2'd0;
wire main_genericstandalone_interface1_bus_err;
reg main_rtio_analyzer_enable_storage_full = 1'd0;
wire main_rtio_analyzer_enable_storage;
reg main_rtio_analyzer_enable_re = 1'd0;
reg main_rtio_analyzer_busy_status = 1'd0;
reg main_rtio_analyzer_message_encoder_source_stb = 1'd0;
wire main_rtio_analyzer_message_encoder_source_ack;
reg main_rtio_analyzer_message_encoder_source_eop = 1'd0;
reg [255:0] main_rtio_analyzer_message_encoder_source_payload_data = 256'd0;
reg main_rtio_analyzer_message_encoder_status = 1'd0;
wire main_rtio_analyzer_message_encoder_overflow_reset_re;
wire main_rtio_analyzer_message_encoder_overflow_reset_r;
reg main_rtio_analyzer_message_encoder_overflow_reset_w = 1'd0;
reg main_rtio_analyzer_message_encoder_read_wait_event_r = 1'd0;
reg main_rtio_analyzer_message_encoder_read_done;
reg main_rtio_analyzer_message_encoder_read_overflow;
wire main_rtio_analyzer_message_encoder_input_output_stb;
reg [1:0] main_rtio_analyzer_message_encoder_input_output_message_type;
wire [29:0] main_rtio_analyzer_message_encoder_input_output_channel;
reg [63:0] main_rtio_analyzer_message_encoder_input_output_timestamp;
wire [63:0] main_rtio_analyzer_message_encoder_input_output_rtio_counter;
wire [31:0] main_rtio_analyzer_message_encoder_input_output_address_padding;
reg [63:0] main_rtio_analyzer_message_encoder_input_output_data;
reg main_rtio_analyzer_message_encoder_exception_stb;
wire [1:0] main_rtio_analyzer_message_encoder_exception_message_type;
wire [29:0] main_rtio_analyzer_message_encoder_exception_channel;
reg [63:0] main_rtio_analyzer_message_encoder_exception_padding0 = 64'd0;
wire [63:0] main_rtio_analyzer_message_encoder_exception_rtio_counter;
reg [7:0] main_rtio_analyzer_message_encoder_exception_exception_type;
reg [87:0] main_rtio_analyzer_message_encoder_exception_padding1 = 88'd0;
reg main_rtio_analyzer_message_encoder_just_written = 1'd0;
wire [1:0] main_rtio_analyzer_message_encoder_stopped_message_type;
reg [93:0] main_rtio_analyzer_message_encoder_stopped_padding0 = 94'd0;
wire [63:0] main_rtio_analyzer_message_encoder_stopped_rtio_counter;
reg [95:0] main_rtio_analyzer_message_encoder_stopped_padding1 = 96'd0;
reg main_rtio_analyzer_message_encoder_enable_r = 1'd0;
reg main_rtio_analyzer_message_encoder_stopping = 1'd0;
wire main_rtio_analyzer_fifo_sink_stb;
wire main_rtio_analyzer_fifo_sink_ack;
wire main_rtio_analyzer_fifo_sink_eop;
wire [255:0] main_rtio_analyzer_fifo_sink_payload_data;
wire main_rtio_analyzer_fifo_source_stb;
wire main_rtio_analyzer_fifo_source_ack;
wire main_rtio_analyzer_fifo_source_eop;
wire [255:0] main_rtio_analyzer_fifo_source_payload_data;
wire main_rtio_analyzer_fifo_re;
reg main_rtio_analyzer_fifo_readable = 1'd0;
wire main_rtio_analyzer_fifo_syncfifo_we;
wire main_rtio_analyzer_fifo_syncfifo_writable;
wire main_rtio_analyzer_fifo_syncfifo_re;
wire main_rtio_analyzer_fifo_syncfifo_readable;
wire [256:0] main_rtio_analyzer_fifo_syncfifo_din;
wire [256:0] main_rtio_analyzer_fifo_syncfifo_dout;
reg [7:0] main_rtio_analyzer_fifo_level0 = 8'd0;
reg main_rtio_analyzer_fifo_replace = 1'd0;
reg [6:0] main_rtio_analyzer_fifo_produce = 7'd0;
reg [6:0] main_rtio_analyzer_fifo_consume = 7'd0;
reg [6:0] main_rtio_analyzer_fifo_wrport_adr;
wire [256:0] main_rtio_analyzer_fifo_wrport_dat_r;
wire main_rtio_analyzer_fifo_wrport_we;
wire [256:0] main_rtio_analyzer_fifo_wrport_dat_w;
wire main_rtio_analyzer_fifo_do_read;
wire [6:0] main_rtio_analyzer_fifo_rdport_adr;
wire [256:0] main_rtio_analyzer_fifo_rdport_dat_r;
wire main_rtio_analyzer_fifo_rdport_re;
wire [7:0] main_rtio_analyzer_fifo_level1;
wire [255:0] main_rtio_analyzer_fifo_fifo_in_payload_data;
wire main_rtio_analyzer_fifo_fifo_in_eop;
wire [255:0] main_rtio_analyzer_fifo_fifo_out_payload_data;
wire main_rtio_analyzer_fifo_fifo_out_eop;
wire main_rtio_analyzer_converter_sink_stb;
wire main_rtio_analyzer_converter_sink_ack;
wire main_rtio_analyzer_converter_sink_eop;
wire [255:0] main_rtio_analyzer_converter_sink_payload_data;
wire main_rtio_analyzer_converter_source_stb;
wire main_rtio_analyzer_converter_source_ack;
wire main_rtio_analyzer_converter_source_eop;
reg [127:0] main_rtio_analyzer_converter_source_payload_data;
wire main_rtio_analyzer_converter_source_payload_valid_token_count;
reg main_rtio_analyzer_converter_mux = 1'd0;
wire main_rtio_analyzer_converter_last;
wire main_rtio_analyzer_dma_reset_re;
wire main_rtio_analyzer_dma_reset_r;
reg main_rtio_analyzer_dma_reset_w = 1'd0;
reg [33:0] main_rtio_analyzer_dma_base_address_storage_full = 34'd0;
wire [29:0] main_rtio_analyzer_dma_base_address_storage;
reg main_rtio_analyzer_dma_base_address_re = 1'd0;
reg [33:0] main_rtio_analyzer_dma_last_address_storage_full = 34'd0;
wire [29:0] main_rtio_analyzer_dma_last_address_storage;
reg main_rtio_analyzer_dma_last_address_re = 1'd0;
wire [63:0] main_rtio_analyzer_dma_status;
wire main_rtio_analyzer_dma_sink_stb;
wire main_rtio_analyzer_dma_sink_ack;
wire main_rtio_analyzer_dma_sink_eop;
wire [127:0] main_rtio_analyzer_dma_sink_payload_data;
wire main_rtio_analyzer_dma_sink_payload_valid_token_count;
reg [58:0] main_rtio_analyzer_dma_message_count = 59'd0;
reg main_rtio_analyzer_enable_r = 1'd0;
reg [5:0] builder_minicon_state = 6'd0;
reg [5:0] builder_minicon_next_state;
reg [2:0] builder_fullmemorywe_state = 3'd0;
reg [2:0] builder_fullmemorywe_next_state;
reg [2:0] builder_a7_1000basex_transmitpath_state = 3'd0;
reg [2:0] builder_a7_1000basex_transmitpath_next_state;
reg main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value;
reg main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce;
reg [2:0] builder_a7_1000basex_receivepath_state = 3'd0;
reg [2:0] builder_a7_1000basex_receivepath_next_state;
reg [1:0] builder_a7_1000basex_fsm_state = 2'd0;
reg [1:0] builder_a7_1000basex_fsm_next_state;
reg [1:0] builder_a7_1000basex_gtptxinit_state = 2'd0;
reg [1:0] builder_a7_1000basex_gtptxinit_next_state;
reg [3:0] builder_a7_1000basex_gtprxinit_state = 4'd0;
reg [3:0] builder_a7_1000basex_gtprxinit_next_state;
reg [15:0] main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value;
reg main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce;
reg builder_liteethmacgap_state = 1'd0;
reg builder_liteethmacgap_next_state;
reg [1:0] builder_liteethmacpreambleinserter_state = 2'd0;
reg [1:0] builder_liteethmacpreambleinserter_next_state;
reg builder_liteethmacpreamblechecker_state = 1'd0;
reg builder_liteethmacpreamblechecker_next_state;
reg [1:0] builder_liteethmaccrc32inserter_state = 2'd0;
reg [1:0] builder_liteethmaccrc32inserter_next_state;
reg [1:0] builder_liteethmaccrc32checker_state = 2'd0;
reg [1:0] builder_liteethmaccrc32checker_next_state;
reg builder_liteethmacpaddinginserter_state = 1'd0;
reg builder_liteethmacpaddinginserter_next_state;
reg [1:0] builder_liteethmacsramwriter_state = 2'd0;
reg [1:0] builder_liteethmacsramwriter_next_state;
reg [31:0] main_genericstandalone_writer_errors_status_next_value;
reg main_genericstandalone_writer_errors_status_next_value_ce;
reg [1:0] builder_liteethmacsramreader_state = 2'd0;
reg [1:0] builder_liteethmacsramreader_next_state;
wire [29:0] builder_shared_adr;
wire [31:0] builder_shared_dat_w;
wire [31:0] builder_shared_dat_r;
wire [3:0] builder_shared_sel;
wire builder_shared_cyc;
wire builder_shared_stb;
wire builder_shared_ack;
wire builder_shared_we;
wire [2:0] builder_shared_cti;
wire [1:0] builder_shared_bte;
wire builder_shared_err;
wire [1:0] builder_request;
reg builder_grant = 1'd0;
reg [4:0] builder_slave_sel;
reg [4:0] builder_slave_sel_r = 5'd0;
reg [2:0] builder_spimaster0_state = 3'd0;
reg [2:0] builder_spimaster0_next_state;
reg [2:0] builder_spimaster1_state = 3'd0;
reg [2:0] builder_spimaster1_next_state;
reg [2:0] builder_spimaster2_state = 3'd0;
reg [2:0] builder_spimaster2_next_state;
reg [1:0] builder_clockdomainsrenamer_resetinserter_state = 2'd0;
reg [1:0] builder_clockdomainsrenamer_resetinserter_next_state;
reg [1:0] builder_clockdomainsrenamer_recordconverter_state = 2'd0;
reg [1:0] builder_clockdomainsrenamer_recordconverter_next_state;
reg [2:0] builder_clockdomainsrenamer_crimaster_state = 3'd0;
reg [2:0] builder_clockdomainsrenamer_crimaster_next_state;
reg [2:0] builder_clockdomainsrenamer_fsm_state = 3'd0;
reg [2:0] builder_clockdomainsrenamer_fsm_next_state;
wire [1:0] builder_sdram_cpulevel_arbiter_request;
reg builder_sdram_cpulevel_arbiter_grant = 1'd0;
wire [2:0] builder_sdram_native_arbiter_request;
reg [1:0] builder_sdram_native_arbiter_grant = 2'd0;
wire [29:0] builder_genericstandalone_shared_adr;
wire [31:0] builder_genericstandalone_shared_dat_w;
wire [31:0] builder_genericstandalone_shared_dat_r;
wire [3:0] builder_genericstandalone_shared_sel;
wire builder_genericstandalone_shared_cyc;
wire builder_genericstandalone_shared_stb;
wire builder_genericstandalone_shared_ack;
wire builder_genericstandalone_shared_we;
wire [2:0] builder_genericstandalone_shared_cti;
wire [1:0] builder_genericstandalone_shared_bte;
wire builder_genericstandalone_shared_err;
wire [1:0] builder_genericstandalone_request;
reg builder_genericstandalone_grant = 1'd0;
reg [5:0] builder_genericstandalone_slave_sel;
reg [5:0] builder_genericstandalone_slave_sel_r = 6'd0;
wire [13:0] builder_genericstandalone_interface0_bank_bus_adr;
wire builder_genericstandalone_interface0_bank_bus_we;
wire [7:0] builder_genericstandalone_interface0_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface0_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank0_dly_sel0_re;
wire [1:0] builder_genericstandalone_csrbank0_dly_sel0_r;
wire [1:0] builder_genericstandalone_csrbank0_dly_sel0_w;
wire builder_genericstandalone_csrbank0_sel;
wire [13:0] builder_genericstandalone_interface1_bank_bus_adr;
wire builder_genericstandalone_interface1_bank_bus_we;
wire [7:0] builder_genericstandalone_interface1_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface1_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank1_control0_re;
wire [3:0] builder_genericstandalone_csrbank1_control0_r;
wire [3:0] builder_genericstandalone_csrbank1_control0_w;
wire builder_genericstandalone_csrbank1_pi0_command0_re;
wire [5:0] builder_genericstandalone_csrbank1_pi0_command0_r;
wire [5:0] builder_genericstandalone_csrbank1_pi0_command0_w;
wire builder_genericstandalone_csrbank1_pi0_address1_re;
wire [6:0] builder_genericstandalone_csrbank1_pi0_address1_r;
wire [6:0] builder_genericstandalone_csrbank1_pi0_address1_w;
wire builder_genericstandalone_csrbank1_pi0_address0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_address0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_address0_w;
wire builder_genericstandalone_csrbank1_pi0_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank1_pi0_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank1_pi0_baddress0_w;
wire builder_genericstandalone_csrbank1_pi0_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata3_w;
wire builder_genericstandalone_csrbank1_pi0_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata2_w;
wire builder_genericstandalone_csrbank1_pi0_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata1_w;
wire builder_genericstandalone_csrbank1_pi0_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_wrdata0_w;
wire builder_genericstandalone_csrbank1_pi0_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata3_w;
wire builder_genericstandalone_csrbank1_pi0_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata2_w;
wire builder_genericstandalone_csrbank1_pi0_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata1_w;
wire builder_genericstandalone_csrbank1_pi0_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi0_rddata0_w;
wire builder_genericstandalone_csrbank1_pi1_command0_re;
wire [5:0] builder_genericstandalone_csrbank1_pi1_command0_r;
wire [5:0] builder_genericstandalone_csrbank1_pi1_command0_w;
wire builder_genericstandalone_csrbank1_pi1_address1_re;
wire [6:0] builder_genericstandalone_csrbank1_pi1_address1_r;
wire [6:0] builder_genericstandalone_csrbank1_pi1_address1_w;
wire builder_genericstandalone_csrbank1_pi1_address0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_address0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_address0_w;
wire builder_genericstandalone_csrbank1_pi1_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank1_pi1_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank1_pi1_baddress0_w;
wire builder_genericstandalone_csrbank1_pi1_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata3_w;
wire builder_genericstandalone_csrbank1_pi1_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata2_w;
wire builder_genericstandalone_csrbank1_pi1_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata1_w;
wire builder_genericstandalone_csrbank1_pi1_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_wrdata0_w;
wire builder_genericstandalone_csrbank1_pi1_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata3_w;
wire builder_genericstandalone_csrbank1_pi1_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata2_w;
wire builder_genericstandalone_csrbank1_pi1_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata1_w;
wire builder_genericstandalone_csrbank1_pi1_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi1_rddata0_w;
wire builder_genericstandalone_csrbank1_pi2_command0_re;
wire [5:0] builder_genericstandalone_csrbank1_pi2_command0_r;
wire [5:0] builder_genericstandalone_csrbank1_pi2_command0_w;
wire builder_genericstandalone_csrbank1_pi2_address1_re;
wire [6:0] builder_genericstandalone_csrbank1_pi2_address1_r;
wire [6:0] builder_genericstandalone_csrbank1_pi2_address1_w;
wire builder_genericstandalone_csrbank1_pi2_address0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_address0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_address0_w;
wire builder_genericstandalone_csrbank1_pi2_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank1_pi2_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank1_pi2_baddress0_w;
wire builder_genericstandalone_csrbank1_pi2_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata3_w;
wire builder_genericstandalone_csrbank1_pi2_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata2_w;
wire builder_genericstandalone_csrbank1_pi2_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata1_w;
wire builder_genericstandalone_csrbank1_pi2_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_wrdata0_w;
wire builder_genericstandalone_csrbank1_pi2_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata3_w;
wire builder_genericstandalone_csrbank1_pi2_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata2_w;
wire builder_genericstandalone_csrbank1_pi2_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata1_w;
wire builder_genericstandalone_csrbank1_pi2_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi2_rddata0_w;
wire builder_genericstandalone_csrbank1_pi3_command0_re;
wire [5:0] builder_genericstandalone_csrbank1_pi3_command0_r;
wire [5:0] builder_genericstandalone_csrbank1_pi3_command0_w;
wire builder_genericstandalone_csrbank1_pi3_address1_re;
wire [6:0] builder_genericstandalone_csrbank1_pi3_address1_r;
wire [6:0] builder_genericstandalone_csrbank1_pi3_address1_w;
wire builder_genericstandalone_csrbank1_pi3_address0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_address0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_address0_w;
wire builder_genericstandalone_csrbank1_pi3_baddress0_re;
wire [2:0] builder_genericstandalone_csrbank1_pi3_baddress0_r;
wire [2:0] builder_genericstandalone_csrbank1_pi3_baddress0_w;
wire builder_genericstandalone_csrbank1_pi3_wrdata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata3_w;
wire builder_genericstandalone_csrbank1_pi3_wrdata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata2_w;
wire builder_genericstandalone_csrbank1_pi3_wrdata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata1_w;
wire builder_genericstandalone_csrbank1_pi3_wrdata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_wrdata0_w;
wire builder_genericstandalone_csrbank1_pi3_rddata3_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata3_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata3_w;
wire builder_genericstandalone_csrbank1_pi3_rddata2_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata2_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata2_w;
wire builder_genericstandalone_csrbank1_pi3_rddata1_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata1_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata1_w;
wire builder_genericstandalone_csrbank1_pi3_rddata0_re;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata0_r;
wire [7:0] builder_genericstandalone_csrbank1_pi3_rddata0_w;
wire builder_genericstandalone_csrbank1_sel;
wire [13:0] builder_genericstandalone_interface2_bank_bus_adr;
wire builder_genericstandalone_interface2_bank_bus_we;
wire [7:0] builder_genericstandalone_interface2_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface2_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank2_sram_writer_slot_re;
wire [1:0] builder_genericstandalone_csrbank2_sram_writer_slot_r;
wire [1:0] builder_genericstandalone_csrbank2_sram_writer_slot_w;
wire builder_genericstandalone_csrbank2_sram_writer_length3_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length3_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length3_w;
wire builder_genericstandalone_csrbank2_sram_writer_length2_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length2_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length2_w;
wire builder_genericstandalone_csrbank2_sram_writer_length1_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length1_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length1_w;
wire builder_genericstandalone_csrbank2_sram_writer_length0_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length0_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_length0_w;
wire builder_genericstandalone_csrbank2_sram_writer_errors3_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors3_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors3_w;
wire builder_genericstandalone_csrbank2_sram_writer_errors2_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors2_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors2_w;
wire builder_genericstandalone_csrbank2_sram_writer_errors1_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors1_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors1_w;
wire builder_genericstandalone_csrbank2_sram_writer_errors0_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors0_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_writer_errors0_w;
wire builder_genericstandalone_csrbank2_sram_writer_ev_enable0_re;
wire builder_genericstandalone_csrbank2_sram_writer_ev_enable0_r;
wire builder_genericstandalone_csrbank2_sram_writer_ev_enable0_w;
wire builder_genericstandalone_csrbank2_sram_reader_ready_re;
wire builder_genericstandalone_csrbank2_sram_reader_ready_r;
wire builder_genericstandalone_csrbank2_sram_reader_ready_w;
wire builder_genericstandalone_csrbank2_sram_reader_slot0_re;
wire [1:0] builder_genericstandalone_csrbank2_sram_reader_slot0_r;
wire [1:0] builder_genericstandalone_csrbank2_sram_reader_slot0_w;
wire builder_genericstandalone_csrbank2_sram_reader_length1_re;
wire [2:0] builder_genericstandalone_csrbank2_sram_reader_length1_r;
wire [2:0] builder_genericstandalone_csrbank2_sram_reader_length1_w;
wire builder_genericstandalone_csrbank2_sram_reader_length0_re;
wire [7:0] builder_genericstandalone_csrbank2_sram_reader_length0_r;
wire [7:0] builder_genericstandalone_csrbank2_sram_reader_length0_w;
wire builder_genericstandalone_csrbank2_sram_reader_ev_enable0_re;
wire builder_genericstandalone_csrbank2_sram_reader_ev_enable0_r;
wire builder_genericstandalone_csrbank2_sram_reader_ev_enable0_w;
wire builder_genericstandalone_csrbank2_preamble_errors3_re;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors3_r;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors3_w;
wire builder_genericstandalone_csrbank2_preamble_errors2_re;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors2_r;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors2_w;
wire builder_genericstandalone_csrbank2_preamble_errors1_re;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors1_r;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors1_w;
wire builder_genericstandalone_csrbank2_preamble_errors0_re;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors0_r;
wire [7:0] builder_genericstandalone_csrbank2_preamble_errors0_w;
wire builder_genericstandalone_csrbank2_crc_errors3_re;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors3_r;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors3_w;
wire builder_genericstandalone_csrbank2_crc_errors2_re;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors2_r;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors2_w;
wire builder_genericstandalone_csrbank2_crc_errors1_re;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors1_r;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors1_w;
wire builder_genericstandalone_csrbank2_crc_errors0_re;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors0_r;
wire [7:0] builder_genericstandalone_csrbank2_crc_errors0_w;
wire builder_genericstandalone_csrbank2_sel;
wire [13:0] builder_genericstandalone_interface3_bank_bus_adr;
wire builder_genericstandalone_interface3_bank_bus_we;
wire [7:0] builder_genericstandalone_interface3_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface3_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank3_in_re;
wire [1:0] builder_genericstandalone_csrbank3_in_r;
wire [1:0] builder_genericstandalone_csrbank3_in_w;
wire builder_genericstandalone_csrbank3_out0_re;
wire [1:0] builder_genericstandalone_csrbank3_out0_r;
wire [1:0] builder_genericstandalone_csrbank3_out0_w;
wire builder_genericstandalone_csrbank3_oe0_re;
wire [1:0] builder_genericstandalone_csrbank3_oe0_r;
wire [1:0] builder_genericstandalone_csrbank3_oe0_w;
wire builder_genericstandalone_csrbank3_sel;
wire [13:0] builder_genericstandalone_interface4_bank_bus_adr;
wire builder_genericstandalone_interface4_bank_bus_we;
wire [7:0] builder_genericstandalone_interface4_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface4_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank4_address0_re;
wire [7:0] builder_genericstandalone_csrbank4_address0_r;
wire [7:0] builder_genericstandalone_csrbank4_address0_w;
wire builder_genericstandalone_csrbank4_data_re;
wire [7:0] builder_genericstandalone_csrbank4_data_r;
wire [7:0] builder_genericstandalone_csrbank4_data_w;
wire builder_genericstandalone_csrbank4_sel;
wire [13:0] builder_genericstandalone_interface5_bank_bus_adr;
wire builder_genericstandalone_interface5_bank_bus_we;
wire [7:0] builder_genericstandalone_interface5_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface5_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank5_reset0_re;
wire builder_genericstandalone_csrbank5_reset0_r;
wire builder_genericstandalone_csrbank5_reset0_w;
wire builder_genericstandalone_csrbank5_sel;
wire [13:0] builder_genericstandalone_interface6_bank_bus_adr;
wire builder_genericstandalone_interface6_bank_bus_we;
wire [7:0] builder_genericstandalone_interface6_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface6_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank6_out0_re;
wire builder_genericstandalone_csrbank6_out0_r;
wire builder_genericstandalone_csrbank6_out0_w;
wire builder_genericstandalone_csrbank6_sel;
wire [13:0] builder_genericstandalone_interface7_bank_bus_adr;
wire builder_genericstandalone_interface7_bank_bus_we;
wire [7:0] builder_genericstandalone_interface7_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface7_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank7_enable0_re;
wire builder_genericstandalone_csrbank7_enable0_r;
wire builder_genericstandalone_csrbank7_enable0_w;
wire builder_genericstandalone_csrbank7_busy_re;
wire builder_genericstandalone_csrbank7_busy_r;
wire builder_genericstandalone_csrbank7_busy_w;
wire builder_genericstandalone_csrbank7_message_encoder_overflow_re;
wire builder_genericstandalone_csrbank7_message_encoder_overflow_r;
wire builder_genericstandalone_csrbank7_message_encoder_overflow_w;
wire builder_genericstandalone_csrbank7_dma_base_address4_re;
wire [1:0] builder_genericstandalone_csrbank7_dma_base_address4_r;
wire [1:0] builder_genericstandalone_csrbank7_dma_base_address4_w;
wire builder_genericstandalone_csrbank7_dma_base_address3_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address3_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address3_w;
wire builder_genericstandalone_csrbank7_dma_base_address2_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address2_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address2_w;
wire builder_genericstandalone_csrbank7_dma_base_address1_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address1_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address1_w;
wire builder_genericstandalone_csrbank7_dma_base_address0_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address0_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_base_address0_w;
wire builder_genericstandalone_csrbank7_dma_last_address4_re;
wire [1:0] builder_genericstandalone_csrbank7_dma_last_address4_r;
wire [1:0] builder_genericstandalone_csrbank7_dma_last_address4_w;
wire builder_genericstandalone_csrbank7_dma_last_address3_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address3_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address3_w;
wire builder_genericstandalone_csrbank7_dma_last_address2_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address2_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address2_w;
wire builder_genericstandalone_csrbank7_dma_last_address1_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address1_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address1_w;
wire builder_genericstandalone_csrbank7_dma_last_address0_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address0_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_last_address0_w;
wire builder_genericstandalone_csrbank7_dma_byte_count7_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count7_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count7_w;
wire builder_genericstandalone_csrbank7_dma_byte_count6_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count6_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count6_w;
wire builder_genericstandalone_csrbank7_dma_byte_count5_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count5_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count5_w;
wire builder_genericstandalone_csrbank7_dma_byte_count4_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count4_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count4_w;
wire builder_genericstandalone_csrbank7_dma_byte_count3_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count3_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count3_w;
wire builder_genericstandalone_csrbank7_dma_byte_count2_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count2_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count2_w;
wire builder_genericstandalone_csrbank7_dma_byte_count1_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count1_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count1_w;
wire builder_genericstandalone_csrbank7_dma_byte_count0_re;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count0_r;
wire [7:0] builder_genericstandalone_csrbank7_dma_byte_count0_w;
wire builder_genericstandalone_csrbank7_sel;
wire [13:0] builder_genericstandalone_interface8_bank_bus_adr;
wire builder_genericstandalone_interface8_bank_bus_we;
wire [7:0] builder_genericstandalone_interface8_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface8_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank8_collision_channel1_re;
wire [7:0] builder_genericstandalone_csrbank8_collision_channel1_r;
wire [7:0] builder_genericstandalone_csrbank8_collision_channel1_w;
wire builder_genericstandalone_csrbank8_collision_channel0_re;
wire [7:0] builder_genericstandalone_csrbank8_collision_channel0_r;
wire [7:0] builder_genericstandalone_csrbank8_collision_channel0_w;
wire builder_genericstandalone_csrbank8_busy_channel1_re;
wire [7:0] builder_genericstandalone_csrbank8_busy_channel1_r;
wire [7:0] builder_genericstandalone_csrbank8_busy_channel1_w;
wire builder_genericstandalone_csrbank8_busy_channel0_re;
wire [7:0] builder_genericstandalone_csrbank8_busy_channel0_r;
wire [7:0] builder_genericstandalone_csrbank8_busy_channel0_w;
wire builder_genericstandalone_csrbank8_sequence_error_channel1_re;
wire [7:0] builder_genericstandalone_csrbank8_sequence_error_channel1_r;
wire [7:0] builder_genericstandalone_csrbank8_sequence_error_channel1_w;
wire builder_genericstandalone_csrbank8_sequence_error_channel0_re;
wire [7:0] builder_genericstandalone_csrbank8_sequence_error_channel0_r;
wire [7:0] builder_genericstandalone_csrbank8_sequence_error_channel0_w;
wire builder_genericstandalone_csrbank8_sel;
wire [13:0] builder_genericstandalone_interface9_bank_bus_adr;
wire builder_genericstandalone_interface9_bank_bus_we;
wire [7:0] builder_genericstandalone_interface9_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface9_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank9_pll_reset0_re;
wire builder_genericstandalone_csrbank9_pll_reset0_r;
wire builder_genericstandalone_csrbank9_pll_reset0_w;
wire builder_genericstandalone_csrbank9_pll_locked_re;
wire builder_genericstandalone_csrbank9_pll_locked_r;
wire builder_genericstandalone_csrbank9_pll_locked_w;
wire builder_genericstandalone_csrbank9_sel;
wire [13:0] builder_genericstandalone_interface10_bank_bus_adr;
wire builder_genericstandalone_interface10_bank_bus_we;
wire [7:0] builder_genericstandalone_interface10_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface10_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank10_mon_chan_sel0_re;
wire [5:0] builder_genericstandalone_csrbank10_mon_chan_sel0_r;
wire [5:0] builder_genericstandalone_csrbank10_mon_chan_sel0_w;
wire builder_genericstandalone_csrbank10_mon_probe_sel0_re;
wire builder_genericstandalone_csrbank10_mon_probe_sel0_r;
wire builder_genericstandalone_csrbank10_mon_probe_sel0_w;
wire builder_genericstandalone_csrbank10_mon_value_re;
wire builder_genericstandalone_csrbank10_mon_value_r;
wire builder_genericstandalone_csrbank10_mon_value_w;
wire builder_genericstandalone_csrbank10_inj_chan_sel0_re;
wire [5:0] builder_genericstandalone_csrbank10_inj_chan_sel0_r;
wire [5:0] builder_genericstandalone_csrbank10_inj_chan_sel0_w;
wire builder_genericstandalone_csrbank10_inj_override_sel0_re;
wire [1:0] builder_genericstandalone_csrbank10_inj_override_sel0_r;
wire [1:0] builder_genericstandalone_csrbank10_inj_override_sel0_w;
wire builder_genericstandalone_csrbank10_sel;
wire [13:0] builder_genericstandalone_interface11_bank_bus_adr;
wire builder_genericstandalone_interface11_bank_bus_we;
wire [7:0] builder_genericstandalone_interface11_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface11_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank11_bitbang0_re;
wire [3:0] builder_genericstandalone_csrbank11_bitbang0_r;
wire [3:0] builder_genericstandalone_csrbank11_bitbang0_w;
wire builder_genericstandalone_csrbank11_miso_re;
wire builder_genericstandalone_csrbank11_miso_r;
wire builder_genericstandalone_csrbank11_miso_w;
wire builder_genericstandalone_csrbank11_bitbang_en0_re;
wire builder_genericstandalone_csrbank11_bitbang_en0_r;
wire builder_genericstandalone_csrbank11_bitbang_en0_w;
wire builder_genericstandalone_csrbank11_sel;
wire [13:0] builder_genericstandalone_interface12_bank_bus_adr;
wire builder_genericstandalone_interface12_bank_bus_we;
wire [7:0] builder_genericstandalone_interface12_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface12_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank12_load7_re;
wire [7:0] builder_genericstandalone_csrbank12_load7_r;
wire [7:0] builder_genericstandalone_csrbank12_load7_w;
wire builder_genericstandalone_csrbank12_load6_re;
wire [7:0] builder_genericstandalone_csrbank12_load6_r;
wire [7:0] builder_genericstandalone_csrbank12_load6_w;
wire builder_genericstandalone_csrbank12_load5_re;
wire [7:0] builder_genericstandalone_csrbank12_load5_r;
wire [7:0] builder_genericstandalone_csrbank12_load5_w;
wire builder_genericstandalone_csrbank12_load4_re;
wire [7:0] builder_genericstandalone_csrbank12_load4_r;
wire [7:0] builder_genericstandalone_csrbank12_load4_w;
wire builder_genericstandalone_csrbank12_load3_re;
wire [7:0] builder_genericstandalone_csrbank12_load3_r;
wire [7:0] builder_genericstandalone_csrbank12_load3_w;
wire builder_genericstandalone_csrbank12_load2_re;
wire [7:0] builder_genericstandalone_csrbank12_load2_r;
wire [7:0] builder_genericstandalone_csrbank12_load2_w;
wire builder_genericstandalone_csrbank12_load1_re;
wire [7:0] builder_genericstandalone_csrbank12_load1_r;
wire [7:0] builder_genericstandalone_csrbank12_load1_w;
wire builder_genericstandalone_csrbank12_load0_re;
wire [7:0] builder_genericstandalone_csrbank12_load0_r;
wire [7:0] builder_genericstandalone_csrbank12_load0_w;
wire builder_genericstandalone_csrbank12_reload7_re;
wire [7:0] builder_genericstandalone_csrbank12_reload7_r;
wire [7:0] builder_genericstandalone_csrbank12_reload7_w;
wire builder_genericstandalone_csrbank12_reload6_re;
wire [7:0] builder_genericstandalone_csrbank12_reload6_r;
wire [7:0] builder_genericstandalone_csrbank12_reload6_w;
wire builder_genericstandalone_csrbank12_reload5_re;
wire [7:0] builder_genericstandalone_csrbank12_reload5_r;
wire [7:0] builder_genericstandalone_csrbank12_reload5_w;
wire builder_genericstandalone_csrbank12_reload4_re;
wire [7:0] builder_genericstandalone_csrbank12_reload4_r;
wire [7:0] builder_genericstandalone_csrbank12_reload4_w;
wire builder_genericstandalone_csrbank12_reload3_re;
wire [7:0] builder_genericstandalone_csrbank12_reload3_r;
wire [7:0] builder_genericstandalone_csrbank12_reload3_w;
wire builder_genericstandalone_csrbank12_reload2_re;
wire [7:0] builder_genericstandalone_csrbank12_reload2_r;
wire [7:0] builder_genericstandalone_csrbank12_reload2_w;
wire builder_genericstandalone_csrbank12_reload1_re;
wire [7:0] builder_genericstandalone_csrbank12_reload1_r;
wire [7:0] builder_genericstandalone_csrbank12_reload1_w;
wire builder_genericstandalone_csrbank12_reload0_re;
wire [7:0] builder_genericstandalone_csrbank12_reload0_r;
wire [7:0] builder_genericstandalone_csrbank12_reload0_w;
wire builder_genericstandalone_csrbank12_en0_re;
wire builder_genericstandalone_csrbank12_en0_r;
wire builder_genericstandalone_csrbank12_en0_w;
wire builder_genericstandalone_csrbank12_value7_re;
wire [7:0] builder_genericstandalone_csrbank12_value7_r;
wire [7:0] builder_genericstandalone_csrbank12_value7_w;
wire builder_genericstandalone_csrbank12_value6_re;
wire [7:0] builder_genericstandalone_csrbank12_value6_r;
wire [7:0] builder_genericstandalone_csrbank12_value6_w;
wire builder_genericstandalone_csrbank12_value5_re;
wire [7:0] builder_genericstandalone_csrbank12_value5_r;
wire [7:0] builder_genericstandalone_csrbank12_value5_w;
wire builder_genericstandalone_csrbank12_value4_re;
wire [7:0] builder_genericstandalone_csrbank12_value4_r;
wire [7:0] builder_genericstandalone_csrbank12_value4_w;
wire builder_genericstandalone_csrbank12_value3_re;
wire [7:0] builder_genericstandalone_csrbank12_value3_r;
wire [7:0] builder_genericstandalone_csrbank12_value3_w;
wire builder_genericstandalone_csrbank12_value2_re;
wire [7:0] builder_genericstandalone_csrbank12_value2_r;
wire [7:0] builder_genericstandalone_csrbank12_value2_w;
wire builder_genericstandalone_csrbank12_value1_re;
wire [7:0] builder_genericstandalone_csrbank12_value1_r;
wire [7:0] builder_genericstandalone_csrbank12_value1_w;
wire builder_genericstandalone_csrbank12_value0_re;
wire [7:0] builder_genericstandalone_csrbank12_value0_r;
wire [7:0] builder_genericstandalone_csrbank12_value0_w;
wire builder_genericstandalone_csrbank12_ev_enable0_re;
wire builder_genericstandalone_csrbank12_ev_enable0_r;
wire builder_genericstandalone_csrbank12_ev_enable0_w;
wire builder_genericstandalone_csrbank12_sel;
wire [13:0] builder_genericstandalone_interface13_bank_bus_adr;
wire builder_genericstandalone_interface13_bank_bus_we;
wire [7:0] builder_genericstandalone_interface13_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface13_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank13_enable_null0_re;
wire builder_genericstandalone_csrbank13_enable_null0_r;
wire builder_genericstandalone_csrbank13_enable_null0_w;
wire builder_genericstandalone_csrbank13_enable_prog0_re;
wire builder_genericstandalone_csrbank13_enable_prog0_r;
wire builder_genericstandalone_csrbank13_enable_prog0_w;
wire builder_genericstandalone_csrbank13_prog_address3_re;
wire [5:0] builder_genericstandalone_csrbank13_prog_address3_r;
wire [5:0] builder_genericstandalone_csrbank13_prog_address3_w;
wire builder_genericstandalone_csrbank13_prog_address2_re;
wire [7:0] builder_genericstandalone_csrbank13_prog_address2_r;
wire [7:0] builder_genericstandalone_csrbank13_prog_address2_w;
wire builder_genericstandalone_csrbank13_prog_address1_re;
wire [7:0] builder_genericstandalone_csrbank13_prog_address1_r;
wire [7:0] builder_genericstandalone_csrbank13_prog_address1_w;
wire builder_genericstandalone_csrbank13_prog_address0_re;
wire [7:0] builder_genericstandalone_csrbank13_prog_address0_r;
wire [7:0] builder_genericstandalone_csrbank13_prog_address0_w;
wire builder_genericstandalone_csrbank13_sel;
wire [13:0] builder_genericstandalone_interface14_bank_bus_adr;
wire builder_genericstandalone_interface14_bank_bus_we;
wire [7:0] builder_genericstandalone_interface14_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface14_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank14_txfull_re;
wire builder_genericstandalone_csrbank14_txfull_r;
wire builder_genericstandalone_csrbank14_txfull_w;
wire builder_genericstandalone_csrbank14_rxempty_re;
wire builder_genericstandalone_csrbank14_rxempty_r;
wire builder_genericstandalone_csrbank14_rxempty_w;
wire builder_genericstandalone_csrbank14_ev_enable0_re;
wire [1:0] builder_genericstandalone_csrbank14_ev_enable0_r;
wire [1:0] builder_genericstandalone_csrbank14_ev_enable0_w;
wire builder_genericstandalone_csrbank14_sel;
wire [13:0] builder_genericstandalone_interface15_bank_bus_adr;
wire builder_genericstandalone_interface15_bank_bus_we;
wire [7:0] builder_genericstandalone_interface15_bank_bus_dat_w;
reg [7:0] builder_genericstandalone_interface15_bank_bus_dat_r = 8'd0;
wire builder_genericstandalone_csrbank15_tuning_word3_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word3_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word3_w;
wire builder_genericstandalone_csrbank15_tuning_word2_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word2_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word2_w;
wire builder_genericstandalone_csrbank15_tuning_word1_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word1_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word1_w;
wire builder_genericstandalone_csrbank15_tuning_word0_re;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word0_r;
wire [7:0] builder_genericstandalone_csrbank15_tuning_word0_w;
wire builder_genericstandalone_csrbank15_sel;
reg [29:0] builder_comb_rhs_array_muxed0;
reg [31:0] builder_comb_rhs_array_muxed1;
reg [3:0] builder_comb_rhs_array_muxed2;
reg builder_comb_rhs_array_muxed3;
reg builder_comb_rhs_array_muxed4;
reg builder_comb_rhs_array_muxed5;
reg [2:0] builder_comb_rhs_array_muxed6;
reg [1:0] builder_comb_rhs_array_muxed7;
wire builder_comb_lhs_array_muxed;
reg builder_comb_rhs_array_muxed8;
reg [1:0] builder_comb_rhs_array_muxed9;
reg [1:0] builder_comb_rhs_array_muxed10;
reg [23:0] builder_comb_rhs_array_muxed11;
reg [63:0] builder_comb_rhs_array_muxed12;
reg [511:0] builder_comb_rhs_array_muxed13;
reg [7:0] builder_comb_rhs_array_muxed14;
reg [63:0] builder_comb_rhs_array_muxed15;
reg builder_comb_rhs_array_muxed16;
reg builder_comb_rhs_array_muxed17;
reg builder_comb_rhs_array_muxed18;
reg builder_comb_rhs_array_muxed19;
reg builder_comb_rhs_array_muxed20;
reg builder_comb_rhs_array_muxed21;
reg builder_comb_rhs_array_muxed22;
reg builder_comb_rhs_array_muxed23;
reg builder_comb_rhs_array_muxed24;
reg builder_comb_rhs_array_muxed25;
reg builder_comb_rhs_array_muxed26;
reg builder_comb_rhs_array_muxed27;
reg builder_comb_rhs_array_muxed28;
reg builder_comb_rhs_array_muxed29;
reg builder_comb_rhs_array_muxed30;
reg builder_comb_rhs_array_muxed31;
reg builder_comb_rhs_array_muxed32;
reg builder_comb_rhs_array_muxed33;
reg builder_comb_rhs_array_muxed34;
reg builder_comb_rhs_array_muxed35;
reg builder_comb_rhs_array_muxed36;
reg builder_comb_rhs_array_muxed37;
reg builder_comb_rhs_array_muxed38;
reg builder_comb_rhs_array_muxed39;
reg builder_comb_rhs_array_muxed40;
reg builder_comb_rhs_array_muxed41;
reg builder_comb_rhs_array_muxed42;
reg builder_comb_rhs_array_muxed43;
reg builder_comb_rhs_array_muxed44;
reg builder_comb_rhs_array_muxed45;
reg builder_comb_rhs_array_muxed46;
reg builder_comb_rhs_array_muxed47;
reg builder_comb_rhs_array_muxed48;
reg builder_comb_rhs_array_muxed49;
reg builder_comb_rhs_array_muxed50;
reg builder_comb_rhs_array_muxed51;
reg builder_comb_rhs_array_muxed52;
reg builder_comb_rhs_array_muxed53;
reg [29:0] builder_comb_rhs_array_muxed54;
reg [31:0] builder_comb_rhs_array_muxed55;
reg [3:0] builder_comb_rhs_array_muxed56;
reg builder_comb_rhs_array_muxed57;
reg builder_comb_rhs_array_muxed58;
reg builder_comb_rhs_array_muxed59;
reg [2:0] builder_comb_rhs_array_muxed60;
reg [1:0] builder_comb_rhs_array_muxed61;
reg [29:0] builder_comb_rhs_array_muxed62;
reg [127:0] builder_comb_rhs_array_muxed63;
reg [15:0] builder_comb_rhs_array_muxed64;
reg builder_comb_rhs_array_muxed65;
reg builder_comb_rhs_array_muxed66;
reg builder_comb_rhs_array_muxed67;
reg [2:0] builder_comb_rhs_array_muxed68;
reg [1:0] builder_comb_rhs_array_muxed69;
reg [29:0] builder_comb_rhs_array_muxed70;
reg [31:0] builder_comb_rhs_array_muxed71;
reg [3:0] builder_comb_rhs_array_muxed72;
reg builder_comb_rhs_array_muxed73;
reg builder_comb_rhs_array_muxed74;
reg builder_comb_rhs_array_muxed75;
reg [2:0] builder_comb_rhs_array_muxed76;
reg [1:0] builder_comb_rhs_array_muxed77;
reg [2:0] builder_sync_t_rhs_array_muxed0;
reg [2:0] builder_sync_f_t_array_muxed0;
reg [2:0] builder_sync_f_rhs_array_muxed0;
reg [4:0] builder_sync_rhs_array_muxed0;
reg [5:0] builder_sync_f_rhs_array_muxed1;
reg builder_sync_f_rhs_array_muxed2;
reg builder_sync_f_rhs_array_muxed3;
reg [3:0] builder_sync_rhs_array_muxed1;
reg builder_sync_rhs_array_muxed2;
reg builder_sync_f_rhs_array_muxed4;
reg builder_sync_basiclowerer_array_muxed0;
reg builder_sync_basiclowerer_array_muxed1;
reg builder_sync_basiclowerer_array_muxed2;
reg builder_sync_basiclowerer_array_muxed3;
reg builder_sync_basiclowerer_array_muxed4;
reg builder_sync_basiclowerer_array_muxed5;
reg builder_sync_basiclowerer_array_muxed6;
reg builder_sync_basiclowerer_array_muxed7;
reg [7:0] builder_sync_f_t_array_muxed1;
reg [6:0] builder_sync_f_t_array_muxed2;
reg [7:0] builder_sync_f_t_array_muxed3;
reg [6:0] builder_sync_f_t_array_muxed4;
reg [7:0] builder_sync_f_t_array_muxed5;
reg [6:0] builder_sync_f_t_array_muxed6;
reg [7:0] builder_sync_f_t_array_muxed7;
reg [6:0] builder_sync_f_t_array_muxed8;
reg [7:0] builder_sync_f_t_array_muxed9;
reg [6:0] builder_sync_f_t_array_muxed10;
reg [7:0] builder_sync_f_t_array_muxed11;
reg [6:0] builder_sync_f_t_array_muxed12;
reg [7:0] builder_sync_f_t_array_muxed13;
reg [6:0] builder_sync_f_t_array_muxed14;
reg [7:0] builder_sync_f_t_array_muxed15;
reg [6:0] builder_sync_f_t_array_muxed16;
reg [7:0] builder_sync_f_t_array_muxed17;
reg [6:0] builder_sync_f_t_array_muxed18;
reg [7:0] builder_sync_f_t_array_muxed19;
reg [6:0] builder_sync_f_t_array_muxed20;
reg [7:0] builder_sync_f_t_array_muxed21;
reg [6:0] builder_sync_f_t_array_muxed22;
reg [7:0] builder_sync_f_t_array_muxed23;
reg [6:0] builder_sync_f_t_array_muxed24;
reg [7:0] builder_sync_f_t_array_muxed25;
reg [6:0] builder_sync_f_t_array_muxed26;
reg [7:0] builder_sync_f_t_array_muxed27;
reg [6:0] builder_sync_f_t_array_muxed28;
reg [7:0] builder_sync_f_t_array_muxed29;
reg [6:0] builder_sync_f_t_array_muxed30;
reg [7:0] builder_sync_f_t_array_muxed31;
reg [6:0] builder_sync_f_t_array_muxed32;
reg [7:0] builder_sync_f_t_array_muxed33;
reg [6:0] builder_sync_f_t_array_muxed34;
reg [7:0] builder_sync_f_t_array_muxed35;
reg [6:0] builder_sync_f_t_array_muxed36;
reg [7:0] builder_sync_f_t_array_muxed37;
reg [6:0] builder_sync_f_t_array_muxed38;
reg [7:0] builder_sync_f_t_array_muxed39;
reg [6:0] builder_sync_f_t_array_muxed40;
reg [7:0] builder_sync_f_t_array_muxed41;
reg [6:0] builder_sync_f_t_array_muxed42;
reg [7:0] builder_sync_f_t_array_muxed43;
reg [6:0] builder_sync_f_t_array_muxed44;
reg [7:0] builder_sync_f_t_array_muxed45;
reg [6:0] builder_sync_f_t_array_muxed46;
reg [7:0] builder_sync_f_t_array_muxed47;
reg [6:0] builder_sync_f_t_array_muxed48;
reg [7:0] builder_sync_f_t_array_muxed49;
reg [6:0] builder_sync_f_t_array_muxed50;
reg [7:0] builder_sync_f_t_array_muxed51;
reg [6:0] builder_sync_f_t_array_muxed52;
reg [7:0] builder_sync_f_t_array_muxed53;
reg [6:0] builder_sync_f_t_array_muxed54;
reg [7:0] builder_sync_f_t_array_muxed55;
reg [6:0] builder_sync_f_t_array_muxed56;
reg [7:0] builder_sync_f_t_array_muxed57;
reg [6:0] builder_sync_f_t_array_muxed58;
reg [7:0] builder_sync_f_t_array_muxed59;
reg [6:0] builder_sync_f_t_array_muxed60;
reg [7:0] builder_sync_f_t_array_muxed61;
reg [6:0] builder_sync_f_t_array_muxed62;
reg [60:0] builder_sync_rhs_array_muxed3;
reg [60:0] builder_sync_rhs_array_muxed4;
reg [60:0] builder_sync_t_lhs_array_muxed = 61'd0;
reg [31:0] builder_sync_t_rhs_array_muxed1;
reg [64:0] builder_sync_t_rhs_array_muxed2;
reg [31:0] builder_sync_rhs_array_muxed5;
reg [31:0] builder_sync_t_t_array_muxed0 = 32'd0;
reg [31:0] builder_sync_rhs_array_muxed6;
reg [31:0] builder_sync_t_t_array_muxed1 = 32'd0;
reg builder_sync_t_rhs_array_muxed3;
reg builder_sync_t_rhs_array_muxed4;
reg builder_sync_t_rhs_array_muxed5;
reg builder_sync_t_rhs_array_muxed6;
reg builder_sync_t_rhs_array_muxed7;
reg builder_sync_t_rhs_array_muxed8;
reg builder_sync_t_rhs_array_muxed9;
reg builder_sync_t_rhs_array_muxed10;
reg builder_sync_t_rhs_array_muxed11;
reg builder_sync_t_rhs_array_muxed12;
reg builder_sync_t_rhs_array_muxed13;
reg builder_sync_t_rhs_array_muxed14;
reg builder_sync_t_rhs_array_muxed15;
reg builder_sync_t_rhs_array_muxed16;
reg builder_sync_t_rhs_array_muxed17;
reg builder_sync_t_rhs_array_muxed18;
reg builder_sync_t_rhs_array_muxed19;
reg builder_sync_t_rhs_array_muxed20;
reg builder_sync_t_rhs_array_muxed21;
reg builder_sync_t_rhs_array_muxed22;
reg builder_sync_t_rhs_array_muxed23;
reg builder_sync_t_rhs_array_muxed24;
reg builder_sync_t_rhs_array_muxed25;
reg builder_sync_t_rhs_array_muxed26;
reg builder_sync_t_rhs_array_muxed27;
reg builder_sync_t_rhs_array_muxed28;
reg builder_sync_t_rhs_array_muxed29;
reg builder_sync_t_rhs_array_muxed30;
reg builder_sync_t_rhs_array_muxed31;
reg builder_sync_t_rhs_array_muxed32;
reg builder_sync_t_rhs_array_muxed33;
reg builder_sync_t_rhs_array_muxed34;
reg builder_sync_t_rhs_array_muxed35;
reg builder_sync_t_rhs_array_muxed36;
reg builder_sync_t_rhs_array_muxed37;
reg builder_sync_t_rhs_array_muxed38;
reg builder_sync_t_rhs_array_muxed39;
reg builder_sync_t_rhs_array_muxed40;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl0_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl0;
wire builder_xilinxasyncresetsynchronizerimpl0_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl3_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl3_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl1;
wire builder_xilinxasyncresetsynchronizerimpl1_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl2;
wire builder_xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl4_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl4_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl5_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl5_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl6_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl6_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl7_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl7_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl8_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl9_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl9_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl10_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl10_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl11_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl11_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl12_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl12_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl13_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl13_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl14_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl14_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl3;
wire builder_xilinxasyncresetsynchronizerimpl3_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl15_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl15_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [60:0] builder_xilinxmultiregimpl16_regs0 = 61'd0;
(* async_reg = "true", dont_touch = "true" *) reg [60:0] builder_xilinxmultiregimpl16_regs1 = 61'd0;
wire builder_xilinxasyncresetsynchronizerimpl4_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl5_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl17_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl17_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl18_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl18_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl19_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl19_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl20_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl20_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl21_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl21_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl22_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl22_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl23_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl23_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl24_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl24_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl25_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl25_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl26_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl26_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl27_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl27_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl28_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl28_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl29_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl29_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl30_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl30_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl31_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl31_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl32_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl32_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl33_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl33_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl34_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl34_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl36_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl36_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl37_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl37_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl38_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl38_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl39_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl39_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl40_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl40_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl41_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl41_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl42_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl42_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl43_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl43_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl44_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl44_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl45_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl45_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl46_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl46_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl47_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl47_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl48_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl48_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl49_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl49_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl50_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl50_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl51_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl51_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl52_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl52_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl53_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl53_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl54_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl54_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl55_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl55_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl56_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl56_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl57_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl57_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl58_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl58_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl59_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl59_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl60_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl60_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl61_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl61_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl62_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl62_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl63_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl63_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl64_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl64_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl65_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl65_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl66_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl66_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl67_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl67_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl68_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl68_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl69_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl69_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl70_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl70_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl71_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl71_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl72_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl72_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl73_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl73_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl74_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl74_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl75_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl75_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl76_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl76_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl77_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl77_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl78_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl78_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl79_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl79_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl80_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl80_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl81_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl81_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl82_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl82_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl83_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl83_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl84_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl84_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl85_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl85_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl86_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl86_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl87_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl87_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl88_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl88_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl89_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl89_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl90_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl90_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl91_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl91_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl92_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl92_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl93_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl93_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl94_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl94_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl95_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl95_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl96_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl96_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl97_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl97_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl98_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl98_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl99_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl99_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl100_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl100_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl101_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl101_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl102_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl102_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl103_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl103_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl104_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl104_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl105_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl105_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl106_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl106_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl107_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl107_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl108_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl108_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl109_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl109_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl110_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl110_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl111_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl111_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl112_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl112_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl113_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl113_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl114_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl114_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl115_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl115_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl116_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl116_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl117_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl117_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl118_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl118_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl119_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl119_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl120_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl120_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl121_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl121_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl122_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl122_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl123_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl123_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl124_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl124_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl125_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl125_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl126_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl126_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl127_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl127_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl128_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl128_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl129_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl129_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl130_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl130_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl131_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl131_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl132_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl132_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl133_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl133_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl134_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl134_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl135_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl135_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl136_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl136_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl137_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl137_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl138_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl138_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl139_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl139_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl140_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl140_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl141_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl141_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl142_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl142_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl143_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl143_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl144_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl144_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl145_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl145_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl146_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl146_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl147_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl147_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl148_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl148_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl149_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl149_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl150_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl150_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl151_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl151_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl152_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl152_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl153_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl153_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl154_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl154_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl155_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl155_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl156_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl156_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl157_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl157_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl158_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl158_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl159_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl159_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl160_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl160_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl161_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl161_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl162_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl162_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl163_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl163_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl164_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl164_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl165_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl165_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl166_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl166_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl167_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl167_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl168_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl168_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl169_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl169_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl170_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl170_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl171_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl171_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl172_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl172_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl173_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl173_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl174_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl174_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl175_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl175_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl176_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl176_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl177_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl177_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl178_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl178_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl179_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl179_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl180_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl180_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl181_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl181_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl182_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl182_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl183_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl183_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl184_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl184_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl185_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl185_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl186_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl186_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl187_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl187_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl188_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl188_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl189_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl189_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl190_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl190_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl191_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl191_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl192_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl192_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl193_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl193_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl194_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl194_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl195_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl195_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl196_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl196_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl197_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl197_regs1 = 1'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address = main_genericstandalone_genericstandalone_genericstandalone_master_p0_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address = main_genericstandalone_genericstandalone_genericstandalone_master_p1_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address = main_genericstandalone_genericstandalone_genericstandalone_master_p2_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address = main_genericstandalone_genericstandalone_genericstandalone_master_p3_address;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cs_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask;
assign main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata = main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid = main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cas_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_ras_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_we_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask;
assign main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_en;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata = main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata_valid = main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid;
assign sfp_ctl_rate_select = 1'd0;
assign sfp_ctl_tx_disable = 1'd0;
assign sfp_ctl_led = ((((~sfp_ctl_los) & (~sfp_ctl_tx_fault)) & (~sfp_ctl_mod_present_n)) & main_genericstandalone_pcs_link_up);

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_interrupt <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_irq;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[1] <= main_genericstandalone_genericstandalone_genericstandalone_timer0_irq;
	main_genericstandalone_genericstandalone_genericstandalone_interrupt[2] <= main_genericstandalone_ev_irq;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_adr = main_genericstandalone_genericstandalone_genericstandalone_i_adr_o[31:2];
assign main_genericstandalone_genericstandalone_genericstandalone_dbus_adr = main_genericstandalone_genericstandalone_genericstandalone_d_adr_o[31:2];
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_adr = main_genericstandalone_genericstandalone_genericstandalone_dbus_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_w = main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_sel = main_genericstandalone_genericstandalone_genericstandalone_dbus_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_cyc = main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_stb = main_genericstandalone_genericstandalone_genericstandalone_dbus_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_we = main_genericstandalone_genericstandalone_genericstandalone_dbus_we;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_cti = main_genericstandalone_genericstandalone_genericstandalone_dbus_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_bte = main_genericstandalone_genericstandalone_genericstandalone_dbus_bte;

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_dbus_ack <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_dbus_err <= 1'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_tmpu_error) begin
		main_genericstandalone_genericstandalone_genericstandalone_dbus_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_dbus_err <= (main_genericstandalone_genericstandalone_genericstandalone_tmpu_ack | main_genericstandalone_genericstandalone_genericstandalone_tmpu_err);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_dbus_ack <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_ack;
		main_genericstandalone_genericstandalone_genericstandalone_dbus_err <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_err;
	end
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sram_we <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[0] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[0]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[1] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[1]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[2] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[2]);
	main_genericstandalone_genericstandalone_genericstandalone_sram_we[3] <= (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we) & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel[3]);
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sram_adr = main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr[9:0];
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w = main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status = (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger = (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status = (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger = (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb);

// synthesis translate_off
reg dummy_d_3;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re & main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r[0])) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_3 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_4;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w <= 2'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status;
	main_genericstandalone_genericstandalone_genericstandalone_uart_status_w[1] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status;
// synthesis translate_off
	dummy_d_4 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_5;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re & main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r[1])) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_5 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_6;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w <= 2'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[0] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending;
	main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[1] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending;
// synthesis translate_off
	dummy_d_6 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_irq = ((main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[0] & main_genericstandalone_genericstandalone_genericstandalone_uart_storage[0]) | (main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w[1] & main_genericstandalone_genericstandalone_genericstandalone_uart_storage[1]));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_status = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_status = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din = {main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data};
assign {main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data} = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_in_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_sink_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_fifo_out_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_7;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= 4'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_7 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_din;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable | main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_re);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_dout = main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level != 5'd16);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_readable = (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din = {main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data};
assign {main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop, main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data} = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_ack = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_in_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_sink_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_stb = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_eop = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_eop;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_payload_data = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_fifo_out_payload_data;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_8;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= 4'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_8 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_din;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable | main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_re);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_dout = main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level != 5'd16);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_readable = (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger = (main_genericstandalone_genericstandalone_genericstandalone_timer0_value != 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status;

// synthesis translate_off
reg dummy_d_9;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re & main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r)) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_9 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending;
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_irq = (main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w & main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage);
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_status = main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
assign main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg = (~main_genericstandalone_genericstandalone_mmcm_locked);
assign main_genericstandalone_genericstandalone_ddrphy_oe = ((main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[1] | main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[2]) | main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[3]);

// synthesis translate_off
reg dummy_d_10;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= 15'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= 3'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= 32'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= 4'd0;
	main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= 1'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_storage[0]) begin
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p0_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p1_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p2_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_slave_p3_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p0_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p1_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p2_rddata_valid;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_bank <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cas_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cs_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_ras_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_we_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_cke <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_odt <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_reset_n <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_wrdata_mask <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask;
		main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_en <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid <= main_genericstandalone_genericstandalone_genericstandalone_master_p3_rddata_valid;
	end
// synthesis translate_off
	dummy_d_10 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cke = main_genericstandalone_genericstandalone_genericstandalone_storage[1];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_odt = main_genericstandalone_genericstandalone_genericstandalone_storage[2];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_reset_n = main_genericstandalone_genericstandalone_genericstandalone_storage[3];

// synthesis translate_off
reg dummy_d_11;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p0_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_11 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p0_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_12;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p1_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_12 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p1_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_13;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p2_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_13 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p2_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_14;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= 1'd1;
	if (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[0]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[1]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[2]);
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= (~main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[3]);
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_we_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_cas_n <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_inti_p3_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_14 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_address = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[4]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_en = (main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re & main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage[5]);
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage;
assign main_genericstandalone_genericstandalone_genericstandalone_inti_p3_wrdata_mask = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0 = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];

// synthesis translate_off
reg dummy_d_15;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6 <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7 <= 1'd0;
	case (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7])
		1'd0: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0 <= 1'd1;
		end
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1 <= 1'd1;
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2 <= 1'd1;
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3 <= 1'd1;
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4 <= 1'd1;
		end
		3'd5: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5 <= 1'd1;
		end
		3'd6: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6 <= 1'd1;
		end
		3'd7: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_15 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit = ((((((((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle = ((((((((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6)) | (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_wait = (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_wait = (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_16;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_address <= {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_16 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_17;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_address <= {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_17 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_18;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_address <= {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_18 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_reset_n = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_odt = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cke = 1'd1;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_cs_n = 1'd0;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_bank = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_19;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= 15'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= 11'd1024;
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[24:10];
		end else begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write | main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read)) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_address <= {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_19 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r = {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_rddata};
assign {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata} = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w;
assign {main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p3_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_wrdata_mask, main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_wrdata_mask} = (~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_hit = ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle) & (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0 == main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1));
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_done = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count == 1'd0);
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_done = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count == 1'd0);

// synthesis translate_off
reg dummy_d_20;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n <= 1'd1;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read <= 1'd0;
	builder_minicon_next_state <= 6'd0;
	builder_minicon_next_state <= builder_minicon_state;
	case (builder_minicon_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_read <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_en <= 1'd1;
			builder_minicon_next_state <= 2'd2;
		end
		2'd2: begin
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_rddata_valid) begin
				main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd1;
				builder_minicon_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_ras_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_we_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p2_wrdata_en <= 1'd1;
			builder_minicon_next_state <= 4'd9;
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack <= 1'd1;
			builder_minicon_next_state <= 1'd0;
		end
		3'd5: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_precharge_all <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd0;
			builder_minicon_next_state <= 4'd14;
		end
		3'd6: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd0;
			builder_minicon_next_state <= 4'd10;
		end
		3'd7: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_activate <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p0_we_n <= 1'd1;
			builder_minicon_next_state <= 4'd12;
		end
		4'd8: begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_ras_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_cas_n <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_dfi_p1_we_n <= 1'd1;
			builder_minicon_next_state <= 5'd16;
		end
		4'd9: begin
			builder_minicon_next_state <= 3'd4;
		end
		4'd10: begin
			builder_minicon_next_state <= 4'd11;
		end
		4'd11: begin
			builder_minicon_next_state <= 3'd7;
		end
		4'd12: begin
			builder_minicon_next_state <= 4'd13;
		end
		4'd13: begin
			builder_minicon_next_state <= 1'd0;
		end
		4'd14: begin
			builder_minicon_next_state <= 4'd15;
		end
		4'd15: begin
			builder_minicon_next_state <= 4'd8;
		end
		5'd16: begin
			builder_minicon_next_state <= 5'd17;
		end
		5'd17: begin
			builder_minicon_next_state <= 5'd18;
		end
		5'd18: begin
			builder_minicon_next_state <= 5'd19;
		end
		5'd19: begin
			builder_minicon_next_state <= 5'd20;
		end
		5'd20: begin
			builder_minicon_next_state <= 5'd21;
		end
		5'd21: begin
			builder_minicon_next_state <= 5'd22;
		end
		5'd22: begin
			builder_minicon_next_state <= 5'd23;
		end
		5'd23: begin
			builder_minicon_next_state <= 5'd24;
		end
		5'd24: begin
			builder_minicon_next_state <= 5'd25;
		end
		5'd25: begin
			builder_minicon_next_state <= 5'd26;
		end
		5'd26: begin
			builder_minicon_next_state <= 5'd27;
		end
		5'd27: begin
			builder_minicon_next_state <= 5'd28;
		end
		5'd28: begin
			builder_minicon_next_state <= 5'd29;
		end
		5'd29: begin
			builder_minicon_next_state <= 5'd30;
		end
		5'd30: begin
			builder_minicon_next_state <= 5'd31;
		end
		5'd31: begin
			builder_minicon_next_state <= 6'd32;
		end
		6'd32: begin
			builder_minicon_next_state <= 6'd33;
		end
		6'd33: begin
			builder_minicon_next_state <= 6'd34;
		end
		6'd34: begin
			builder_minicon_next_state <= 6'd35;
		end
		6'd35: begin
			builder_minicon_next_state <= 6'd36;
		end
		6'd36: begin
			builder_minicon_next_state <= 6'd37;
		end
		6'd37: begin
			builder_minicon_next_state <= 6'd38;
		end
		6'd38: begin
			builder_minicon_next_state <= 6'd39;
		end
		6'd39: begin
			builder_minicon_next_state <= 6'd40;
		end
		6'd40: begin
			builder_minicon_next_state <= 6'd41;
		end
		6'd41: begin
			builder_minicon_next_state <= 6'd42;
		end
		6'd42: begin
			builder_minicon_next_state <= 6'd43;
		end
		6'd43: begin
			builder_minicon_next_state <= 6'd44;
		end
		6'd44: begin
			builder_minicon_next_state <= 6'd45;
		end
		6'd45: begin
			builder_minicon_next_state <= 1'd0;
		end
		default: begin
			if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_done) begin
				builder_minicon_next_state <= 3'd5;
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb & main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc)) begin
					if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_hit) begin
						if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we) begin
							builder_minicon_next_state <= 2'd3;
						end else begin
							builder_minicon_next_state <= 1'd1;
						end
					end else begin
						if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank_idle)) begin
							if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_done) begin
								builder_minicon_next_state <= 3'd6;
							end
						end else begin
							builder_minicon_next_state <= 3'd7;
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_20 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_data_port_adr = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[14:2];

// synthesis translate_off
reg dummy_d_21;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_data_port_we <= 16'd0;
	main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w <= 128'd0;
	if (main_genericstandalone_genericstandalone_genericstandalone_write_from_slave) begin
		main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r;
		main_genericstandalone_genericstandalone_genericstandalone_data_port_we <= {16{1'd1}};
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w <= {4{main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w}};
		if ((((main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb) & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we) & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack)) begin
			main_genericstandalone_genericstandalone_genericstandalone_data_port_we <= {({4{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[1:0] == 1'd0)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({4{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[1:0] == 1'd1)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({4{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[1:0] == 2'd2)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel), ({4{(main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[1:0] == 2'd3)}} & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel)};
		end
	end
// synthesis translate_off
	dummy_d_21 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel = 16'd65535;

// synthesis translate_off
reg dummy_d_22;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= 32'd0;
	case (main_genericstandalone_genericstandalone_genericstandalone_adr_offset_r)
		1'd0: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[127:96];
		end
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[95:64];
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[63:32];
		end
		default: begin
			main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[31:0];
		end
	endcase
// synthesis translate_off
	dummy_d_22 <= dummy_s;
// synthesis translate_on
end
assign {main_genericstandalone_genericstandalone_genericstandalone_tag_do_dirty, main_genericstandalone_genericstandalone_genericstandalone_tag_do_tag} = main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_w = {main_genericstandalone_genericstandalone_genericstandalone_tag_di_dirty, main_genericstandalone_genericstandalone_genericstandalone_tag_di_tag};
assign main_genericstandalone_genericstandalone_genericstandalone_tag_port_adr = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[14:2];
assign main_genericstandalone_genericstandalone_genericstandalone_tag_di_tag = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[29:15];
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr = {main_genericstandalone_genericstandalone_genericstandalone_tag_do_tag, main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[14:2]};

// synthesis translate_off
reg dummy_d_23;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_write_from_slave <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_tag_port_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_tag_di_dirty <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_word_clr <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_word_inc <= 1'd0;
	builder_fullmemorywe_next_state <= 3'd0;
	builder_fullmemorywe_next_state <= builder_fullmemorywe_state;
	case (builder_fullmemorywe_state)
		1'd1: begin
			main_genericstandalone_genericstandalone_genericstandalone_word_clr <= 1'd1;
			if ((main_genericstandalone_genericstandalone_genericstandalone_tag_do_tag == main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[29:15])) begin
				main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack <= 1'd1;
				if (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we) begin
					main_genericstandalone_genericstandalone_genericstandalone_tag_di_dirty <= 1'd1;
					main_genericstandalone_genericstandalone_genericstandalone_tag_port_we <= 1'd1;
				end
				builder_fullmemorywe_next_state <= 1'd0;
			end else begin
				if (main_genericstandalone_genericstandalone_genericstandalone_tag_do_dirty) begin
					builder_fullmemorywe_next_state <= 2'd2;
				end else begin
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd1;
			if (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack) begin
				main_genericstandalone_genericstandalone_genericstandalone_word_inc <= 1'd1;
				if (1'd1) begin
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			main_genericstandalone_genericstandalone_genericstandalone_tag_port_we <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_word_clr <= 1'd1;
			builder_fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we <= 1'd0;
			if (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack) begin
				main_genericstandalone_genericstandalone_genericstandalone_write_from_slave <= 1'd1;
				main_genericstandalone_genericstandalone_genericstandalone_word_inc <= 1'd1;
				if (1'd1) begin
					builder_fullmemorywe_next_state <= 1'd1;
				end else begin
					builder_fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc & main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb)) begin
				builder_fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_23 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_spiflash_bus_dat_r = main_genericstandalone_genericstandalone_spiflash_sr;

// synthesis translate_off
reg dummy_d_24;
// synthesis translate_on
always @(*) begin
	spiflash2x_cs_n <= 1'd1;
	main_genericstandalone_genericstandalone_clk <= 1'd0;
	main_genericstandalone_genericstandalone_spiflash_status <= 1'd0;
	main_genericstandalone_genericstandalone_spiflash_o <= 2'd0;
	main_genericstandalone_genericstandalone_spiflash_oe <= 1'd0;
	if (main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage) begin
		main_genericstandalone_genericstandalone_clk <= main_genericstandalone_genericstandalone_spiflash_bitbang_storage[1];
		spiflash2x_cs_n <= main_genericstandalone_genericstandalone_spiflash_bitbang_storage[2];
		if (main_genericstandalone_genericstandalone_spiflash_bitbang_storage[3]) begin
			main_genericstandalone_genericstandalone_spiflash_oe <= 1'd0;
		end else begin
			main_genericstandalone_genericstandalone_spiflash_oe <= 1'd1;
		end
		if (main_genericstandalone_genericstandalone_spiflash_bitbang_storage[1]) begin
			main_genericstandalone_genericstandalone_spiflash_status <= main_genericstandalone_genericstandalone_spiflash_i0[1];
		end
		main_genericstandalone_genericstandalone_spiflash_o <= {{1{1'd1}}, main_genericstandalone_genericstandalone_spiflash_bitbang_storage[0]};
	end else begin
		main_genericstandalone_genericstandalone_clk <= main_genericstandalone_genericstandalone_spiflash_clk;
		spiflash2x_cs_n <= main_genericstandalone_genericstandalone_spiflash_cs_n;
		main_genericstandalone_genericstandalone_spiflash_o <= main_genericstandalone_genericstandalone_spiflash_sr[31:30];
		main_genericstandalone_genericstandalone_spiflash_oe <= main_genericstandalone_genericstandalone_spiflash_dq_oe;
	end
// synthesis translate_off
	dummy_d_24 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_qpll_reset = main_genericstandalone_tx_init_qpll_reset0;
assign main_genericstandalone_tx_init_qpll_lock0 = main_genericstandalone_genericstandalone_qpll_lock;
assign main_genericstandalone_tx_reset = main_genericstandalone_tx_init_tx_reset0;
assign main_genericstandalone_rx_init_enable = main_genericstandalone_tx_init_done;
assign main_genericstandalone_rx_reset = main_genericstandalone_rx_init_rx_reset0;
assign main_genericstandalone_rx_init_rx_pma_reset_done0 = main_genericstandalone_rx_pma_reset_done;
assign main_genericstandalone_drpaddr = main_genericstandalone_rx_init_drpaddr;
assign main_genericstandalone_drpen = main_genericstandalone_rx_init_drpen;
assign main_genericstandalone_drpdi = main_genericstandalone_rx_init_drpdi;
assign main_genericstandalone_rx_init_drprdy = main_genericstandalone_drprdy;
assign main_genericstandalone_rx_init_drpdo = main_genericstandalone_drpdo;
assign main_genericstandalone_drpwe = main_genericstandalone_rx_init_drpwe;
assign main_genericstandalone_i = main_genericstandalone_pcs_restart;
assign main_genericstandalone_rx_init_restart = main_genericstandalone_o;
assign main_genericstandalone_tx_data0 = main_genericstandalone_tx_data_half;
assign main_genericstandalone_rx_data_half = main_genericstandalone_rx_data0;
assign main_genericstandalone_tx_data1 = main_genericstandalone_pcs_transmitpath_output0;
assign main_genericstandalone_pcs_receivepath_input = main_genericstandalone_rx_data1;
assign main_genericstandalone_pcs_transmitpath_tx_stb = main_genericstandalone_pcs_sink_stb;
assign main_genericstandalone_pcs_sink_ack = main_genericstandalone_pcs_transmitpath_tx_ack;
assign main_genericstandalone_pcs_transmitpath_tx_data = main_genericstandalone_pcs_sink_payload_data;
assign main_genericstandalone_pcs_source_eop = ((~main_genericstandalone_pcs_receivepath_rx_en) & main_genericstandalone_pcs_rx_en_d);
assign main_genericstandalone_pcs_seen_valid_ci_i = main_genericstandalone_pcs_receivepath_seen_valid_ci;
assign main_genericstandalone_pcs_transmitpath_config_reg = (6'd32 | (main_genericstandalone_pcs_autoneg_ack <<< 4'd14));
assign main_genericstandalone_pcs_transmitpath_d1 = main_genericstandalone_pcs_transmitpath_d0;
assign main_genericstandalone_pcs_transmitpath_k1 = main_genericstandalone_pcs_transmitpath_k0;
assign main_genericstandalone_pcs_transmitpath_disp_inter = (main_genericstandalone_pcs_transmitpath_disp_in ^ main_genericstandalone_pcs_transmitpath_code6b_unbalanced);

// synthesis translate_off
reg dummy_d_25;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_output_6b <= 6'd0;
	if (((~main_genericstandalone_pcs_transmitpath_disp_in) & main_genericstandalone_pcs_transmitpath_code6b_flip)) begin
		main_genericstandalone_pcs_transmitpath_output_6b <= (~main_genericstandalone_pcs_transmitpath_code6b);
	end else begin
		main_genericstandalone_pcs_transmitpath_output_6b <= main_genericstandalone_pcs_transmitpath_code6b;
	end
// synthesis translate_off
	dummy_d_25 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_26;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_disp_out <= 1'd0;
	main_genericstandalone_pcs_transmitpath_output_4b <= 4'd0;
	if (((~main_genericstandalone_pcs_transmitpath_disp_inter) & main_genericstandalone_pcs_transmitpath_alt7_rd0)) begin
		main_genericstandalone_pcs_transmitpath_disp_out <= (~main_genericstandalone_pcs_transmitpath_disp_inter);
		main_genericstandalone_pcs_transmitpath_output_4b <= 3'd7;
	end else begin
		if ((main_genericstandalone_pcs_transmitpath_disp_inter & main_genericstandalone_pcs_transmitpath_alt7_rd1)) begin
			main_genericstandalone_pcs_transmitpath_disp_out <= (~main_genericstandalone_pcs_transmitpath_disp_inter);
			main_genericstandalone_pcs_transmitpath_output_4b <= 4'd8;
		end else begin
			main_genericstandalone_pcs_transmitpath_disp_out <= (main_genericstandalone_pcs_transmitpath_disp_inter ^ main_genericstandalone_pcs_transmitpath_code4b_unbalanced);
			if (((~main_genericstandalone_pcs_transmitpath_disp_inter) & main_genericstandalone_pcs_transmitpath_code4b_flip)) begin
				main_genericstandalone_pcs_transmitpath_output_4b <= (~main_genericstandalone_pcs_transmitpath_code4b);
			end else begin
				main_genericstandalone_pcs_transmitpath_output_4b <= main_genericstandalone_pcs_transmitpath_code4b;
			end
		end
	end
// synthesis translate_off
	dummy_d_26 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_transmitpath_output_msb_first = {main_genericstandalone_pcs_transmitpath_output_6b, main_genericstandalone_pcs_transmitpath_output_4b};

// synthesis translate_off
reg dummy_d_27;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_output1 <= 10'd0;
	main_genericstandalone_pcs_transmitpath_output1[0] <= main_genericstandalone_pcs_transmitpath_output_msb_first[9];
	main_genericstandalone_pcs_transmitpath_output1[1] <= main_genericstandalone_pcs_transmitpath_output_msb_first[8];
	main_genericstandalone_pcs_transmitpath_output1[2] <= main_genericstandalone_pcs_transmitpath_output_msb_first[7];
	main_genericstandalone_pcs_transmitpath_output1[3] <= main_genericstandalone_pcs_transmitpath_output_msb_first[6];
	main_genericstandalone_pcs_transmitpath_output1[4] <= main_genericstandalone_pcs_transmitpath_output_msb_first[5];
	main_genericstandalone_pcs_transmitpath_output1[5] <= main_genericstandalone_pcs_transmitpath_output_msb_first[4];
	main_genericstandalone_pcs_transmitpath_output1[6] <= main_genericstandalone_pcs_transmitpath_output_msb_first[3];
	main_genericstandalone_pcs_transmitpath_output1[7] <= main_genericstandalone_pcs_transmitpath_output_msb_first[2];
	main_genericstandalone_pcs_transmitpath_output1[8] <= main_genericstandalone_pcs_transmitpath_output_msb_first[1];
	main_genericstandalone_pcs_transmitpath_output1[9] <= main_genericstandalone_pcs_transmitpath_output_msb_first[0];
// synthesis translate_off
	dummy_d_27 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_28;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd0;
	main_genericstandalone_pcs_transmitpath_d0 <= 8'd0;
	main_genericstandalone_pcs_transmitpath_k0 <= 1'd0;
	main_genericstandalone_pcs_transmitpath_load_config_reg_buffer <= 1'd0;
	builder_a7_1000basex_transmitpath_next_state <= 3'd0;
	main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value <= 1'd0;
	main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd0;
	builder_a7_1000basex_transmitpath_next_state <= builder_a7_1000basex_transmitpath_state;
	case (builder_a7_1000basex_transmitpath_state)
		1'd1: begin
			if (main_genericstandalone_pcs_transmitpath_c_type) begin
				main_genericstandalone_pcs_transmitpath_d0 <= 7'd66;
			end else begin
				main_genericstandalone_pcs_transmitpath_d0 <= 8'd181;
			end
			main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value <= (~main_genericstandalone_pcs_transmitpath_c_type);
			main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd1;
			builder_a7_1000basex_transmitpath_next_state <= 2'd2;
		end
		2'd2: begin
			main_genericstandalone_pcs_transmitpath_d0 <= main_genericstandalone_pcs_transmitpath_config_reg_buffer[7:0];
			builder_a7_1000basex_transmitpath_next_state <= 2'd3;
		end
		2'd3: begin
			main_genericstandalone_pcs_transmitpath_d0 <= main_genericstandalone_pcs_transmitpath_config_reg_buffer[15:8];
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd4: begin
			if (main_genericstandalone_pcs_transmitpath_disparity) begin
				main_genericstandalone_pcs_transmitpath_d0 <= 8'd197;
			end else begin
				main_genericstandalone_pcs_transmitpath_d0 <= 7'd80;
			end
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd5: begin
			main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd1;
			if (main_genericstandalone_pcs_transmitpath_tx_stb) begin
				main_genericstandalone_pcs_transmitpath_d0 <= main_genericstandalone_pcs_transmitpath_tx_data;
			end else begin
				main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
				main_genericstandalone_pcs_transmitpath_d0 <= 8'd253;
				builder_a7_1000basex_transmitpath_next_state <= 3'd6;
			end
		end
		3'd6: begin
			main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_d0 <= 8'd247;
			if (main_genericstandalone_pcs_transmitpath_parity) begin
				builder_a7_1000basex_transmitpath_next_state <= 1'd0;
			end else begin
				builder_a7_1000basex_transmitpath_next_state <= 3'd7;
			end
		end
		3'd7: begin
			main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_d0 <= 8'd247;
			builder_a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		default: begin
			main_genericstandalone_pcs_transmitpath_tx_ack <= 1'd1;
			if (main_genericstandalone_pcs_transmitpath_config_stb) begin
				main_genericstandalone_pcs_transmitpath_load_config_reg_buffer <= 1'd1;
				main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
				main_genericstandalone_pcs_transmitpath_d0 <= 8'd188;
				builder_a7_1000basex_transmitpath_next_state <= 1'd1;
			end else begin
				if (main_genericstandalone_pcs_transmitpath_tx_stb) begin
					main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
					main_genericstandalone_pcs_transmitpath_d0 <= 8'd251;
					builder_a7_1000basex_transmitpath_next_state <= 3'd5;
				end else begin
					main_genericstandalone_pcs_transmitpath_k0 <= 1'd1;
					main_genericstandalone_pcs_transmitpath_d0 <= 8'd188;
					builder_a7_1000basex_transmitpath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_28 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_receivepath_rx_data = (main_genericstandalone_pcs_receivepath_first_preamble_byte ? 7'd85 : main_genericstandalone_pcs_receivepath_d);

// synthesis translate_off
reg dummy_d_29;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_receivepath_input_msb_first <= 10'd0;
	main_genericstandalone_pcs_receivepath_input_msb_first[0] <= main_genericstandalone_pcs_receivepath_input[9];
	main_genericstandalone_pcs_receivepath_input_msb_first[1] <= main_genericstandalone_pcs_receivepath_input[8];
	main_genericstandalone_pcs_receivepath_input_msb_first[2] <= main_genericstandalone_pcs_receivepath_input[7];
	main_genericstandalone_pcs_receivepath_input_msb_first[3] <= main_genericstandalone_pcs_receivepath_input[6];
	main_genericstandalone_pcs_receivepath_input_msb_first[4] <= main_genericstandalone_pcs_receivepath_input[5];
	main_genericstandalone_pcs_receivepath_input_msb_first[5] <= main_genericstandalone_pcs_receivepath_input[4];
	main_genericstandalone_pcs_receivepath_input_msb_first[6] <= main_genericstandalone_pcs_receivepath_input[3];
	main_genericstandalone_pcs_receivepath_input_msb_first[7] <= main_genericstandalone_pcs_receivepath_input[2];
	main_genericstandalone_pcs_receivepath_input_msb_first[8] <= main_genericstandalone_pcs_receivepath_input[1];
	main_genericstandalone_pcs_receivepath_input_msb_first[9] <= main_genericstandalone_pcs_receivepath_input[0];
// synthesis translate_off
	dummy_d_29 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_receivepath_d = {main_genericstandalone_pcs_receivepath_code3b, main_genericstandalone_pcs_receivepath_code5b};

// synthesis translate_off
reg dummy_d_30;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_receivepath_rx_en <= 1'd0;
	main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd0;
	main_genericstandalone_pcs_receivepath_load_config_reg_lsb <= 1'd0;
	main_genericstandalone_pcs_receivepath_load_config_reg_msb <= 1'd0;
	main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd0;
	builder_a7_1000basex_receivepath_next_state <= 3'd0;
	builder_a7_1000basex_receivepath_next_state <= builder_a7_1000basex_receivepath_state;
	case (builder_a7_1000basex_receivepath_state)
		1'd1: begin
			builder_a7_1000basex_receivepath_next_state <= 1'd0;
			if ((~main_genericstandalone_pcs_receivepath_k)) begin
				if (((main_genericstandalone_pcs_receivepath_d == 8'd181) | (main_genericstandalone_pcs_receivepath_d == 7'd66))) begin
					main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 2'd2;
				end
				if (((main_genericstandalone_pcs_receivepath_d == 8'd197) | (main_genericstandalone_pcs_receivepath_d == 7'd80))) begin
					main_genericstandalone_pcs_receivepath_seen_valid_ci <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end
		end
		2'd2: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				if ((main_genericstandalone_pcs_receivepath_d == 8'd251)) begin
					main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 3'd4;
				end else begin
					builder_a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end else begin
				main_genericstandalone_pcs_receivepath_load_config_reg_lsb <= 1'd1;
				builder_a7_1000basex_receivepath_next_state <= 2'd3;
			end
		end
		2'd3: begin
			if ((~main_genericstandalone_pcs_receivepath_k)) begin
				main_genericstandalone_pcs_receivepath_load_config_reg_msb <= 1'd1;
			end
			builder_a7_1000basex_receivepath_next_state <= 1'd0;
		end
		3'd4: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				builder_a7_1000basex_receivepath_next_state <= 1'd0;
			end else begin
				main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
			end
		end
		default: begin
			if (main_genericstandalone_pcs_receivepath_k) begin
				if ((main_genericstandalone_pcs_receivepath_d == 8'd188)) begin
					builder_a7_1000basex_receivepath_next_state <= 1'd1;
				end
				if ((main_genericstandalone_pcs_receivepath_d == 8'd251)) begin
					main_genericstandalone_pcs_receivepath_rx_en <= 1'd1;
					main_genericstandalone_pcs_receivepath_first_preamble_byte <= 1'd1;
					builder_a7_1000basex_receivepath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_30 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_pcs_seen_valid_ci_o = (main_genericstandalone_pcs_seen_valid_ci_toggle_o ^ main_genericstandalone_pcs_seen_valid_ci_toggle_o_r);
assign main_genericstandalone_pcs_rx_config_reg_o = (main_genericstandalone_pcs_rx_config_reg_toggle_o ^ main_genericstandalone_pcs_rx_config_reg_toggle_o_r);
assign main_genericstandalone_pcs_rx_config_reg_ack_o = (main_genericstandalone_pcs_rx_config_reg_ack_toggle_o ^ main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r);
assign main_genericstandalone_pcs_done = (main_genericstandalone_pcs_count == 1'd0);

// synthesis translate_off
reg dummy_d_31;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_pcs_transmitpath_config_stb <= 1'd0;
	main_genericstandalone_pcs_link_up <= 1'd0;
	main_genericstandalone_pcs_restart <= 1'd0;
	main_genericstandalone_pcs_autoneg_ack <= 1'd0;
	main_genericstandalone_pcs_wait <= 1'd0;
	builder_a7_1000basex_fsm_next_state <= 2'd0;
	builder_a7_1000basex_fsm_next_state <= builder_a7_1000basex_fsm_state;
	case (builder_a7_1000basex_fsm_state)
		1'd1: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			main_genericstandalone_pcs_autoneg_ack <= 1'd1;
			if (main_genericstandalone_pcs_rx_config_reg_ack_o) begin
				builder_a7_1000basex_fsm_next_state <= 2'd2;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd2: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			main_genericstandalone_pcs_autoneg_ack <= 1'd1;
			main_genericstandalone_pcs_wait <= 1'd1;
			if (main_genericstandalone_pcs_done) begin
				builder_a7_1000basex_fsm_next_state <= 2'd3;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_pcs_link_up <= 1'd1;
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_pcs_transmitpath_config_stb <= 1'd1;
			if ((main_genericstandalone_pcs_rx_config_reg_o | main_genericstandalone_pcs_rx_config_reg_ack_o)) begin
				builder_a7_1000basex_fsm_next_state <= 1'd1;
			end
			if ((main_genericstandalone_pcs_checker_tick & (~main_genericstandalone_pcs_checker_ok))) begin
				main_genericstandalone_pcs_restart <= 1'd1;
				builder_a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_31 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_32;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_init_done <= 1'd0;
	main_genericstandalone_tx_init_qpll_reset1 <= 1'd0;
	main_genericstandalone_tx_init_tx_reset1 <= 1'd0;
	builder_a7_1000basex_gtptxinit_next_state <= 2'd0;
	builder_a7_1000basex_gtptxinit_next_state <= builder_a7_1000basex_gtptxinit_state;
	case (builder_a7_1000basex_gtptxinit_state)
		1'd1: begin
			main_genericstandalone_tx_init_tx_reset1 <= 1'd1;
			main_genericstandalone_tx_init_qpll_reset1 <= 1'd1;
			if (main_genericstandalone_tx_init_tick) begin
				builder_a7_1000basex_gtptxinit_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_tx_init_tx_reset1 <= 1'd1;
			if ((main_genericstandalone_tx_init_qpll_lock1 & main_genericstandalone_tx_init_tick)) begin
				builder_a7_1000basex_gtptxinit_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_genericstandalone_tx_init_done <= 1'd1;
		end
		default: begin
			if (main_genericstandalone_tx_init_tick) begin
				builder_a7_1000basex_gtptxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_32 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_init_drpaddr = 5'd17;

// synthesis translate_off
reg dummy_d_33;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_init_drpdi <= 16'd0;
	if (main_genericstandalone_rx_init_drpmask) begin
		main_genericstandalone_rx_init_drpdi <= (main_genericstandalone_rx_init_drpvalue & 16'd63487);
	end else begin
		main_genericstandalone_rx_init_drpdi <= main_genericstandalone_rx_init_drpvalue;
	end
// synthesis translate_off
	dummy_d_33 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_34;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_init_drpen <= 1'd0;
	main_genericstandalone_rx_init_drpwe <= 1'd0;
	main_genericstandalone_rx_init_done <= 1'd0;
	main_genericstandalone_rx_init_rx_reset1 <= 1'd0;
	main_genericstandalone_rx_init_drpmask <= 1'd0;
	builder_a7_1000basex_gtprxinit_next_state <= 4'd0;
	main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value <= 16'd0;
	main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd0;
	builder_a7_1000basex_gtprxinit_next_state <= builder_a7_1000basex_gtprxinit_state;
	case (builder_a7_1000basex_gtprxinit_state)
		1'd1: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 2'd2;
		end
		2'd2: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			main_genericstandalone_rx_init_drpen <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 2'd3;
		end
		2'd3: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			if (main_genericstandalone_rx_init_drprdy) begin
				main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value <= main_genericstandalone_rx_init_drpdo;
				main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd1;
				builder_a7_1000basex_gtprxinit_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			main_genericstandalone_rx_init_drpmask <= 1'd1;
			main_genericstandalone_rx_init_drpen <= 1'd1;
			main_genericstandalone_rx_init_drpwe <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 3'd5;
		end
		3'd5: begin
			main_genericstandalone_rx_init_rx_reset1 <= 1'd1;
			if (main_genericstandalone_rx_init_drprdy) begin
				builder_a7_1000basex_gtprxinit_next_state <= 3'd6;
			end
		end
		3'd6: begin
			if ((main_genericstandalone_rx_init_rx_pma_reset_done_r & (~main_genericstandalone_rx_init_rx_pma_reset_done1))) begin
				builder_a7_1000basex_gtprxinit_next_state <= 3'd7;
			end
		end
		3'd7: begin
			main_genericstandalone_rx_init_drpen <= 1'd1;
			main_genericstandalone_rx_init_drpwe <= 1'd1;
			builder_a7_1000basex_gtprxinit_next_state <= 4'd8;
		end
		4'd8: begin
			if (main_genericstandalone_rx_init_drprdy) begin
				builder_a7_1000basex_gtprxinit_next_state <= 4'd9;
			end
		end
		4'd9: begin
			main_genericstandalone_rx_init_done <= 1'd1;
			if (main_genericstandalone_rx_init_restart) begin
				builder_a7_1000basex_gtprxinit_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_genericstandalone_rx_init_enable) begin
				builder_a7_1000basex_gtprxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_34 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_o = (main_genericstandalone_toggle_o ^ main_genericstandalone_toggle_o_r);
assign main_genericstandalone_tx_cdc_sink_stb = main_genericstandalone_source_stb;
assign main_genericstandalone_source_ack = main_genericstandalone_tx_cdc_sink_ack;
assign main_genericstandalone_tx_cdc_sink_eop = main_genericstandalone_source_eop;
assign main_genericstandalone_tx_cdc_sink_payload_data = main_genericstandalone_source_payload_data;
assign main_genericstandalone_tx_cdc_sink_payload_last_be = main_genericstandalone_source_payload_last_be;
assign main_genericstandalone_tx_cdc_sink_payload_error = main_genericstandalone_source_payload_error;
assign main_genericstandalone_sink_stb = main_genericstandalone_rx_cdc_source_stb;
assign main_genericstandalone_rx_cdc_source_ack = main_genericstandalone_sink_ack;
assign main_genericstandalone_sink_eop = main_genericstandalone_rx_cdc_source_eop;
assign main_genericstandalone_sink_payload_data = main_genericstandalone_rx_cdc_source_payload_data;
assign main_genericstandalone_sink_payload_last_be = main_genericstandalone_rx_cdc_source_payload_last_be;
assign main_genericstandalone_sink_payload_error = main_genericstandalone_rx_cdc_source_payload_error;
assign main_genericstandalone_ps_preamble_error_i = main_genericstandalone_preamble_checker_error;
assign main_genericstandalone_ps_crc_error_i = main_genericstandalone_crc32_checker_error;
assign main_genericstandalone_tx_converter_sink_sink_stb = main_genericstandalone_tx_cdc_source_stb;
assign main_genericstandalone_tx_cdc_source_ack = main_genericstandalone_tx_converter_sink_sink_ack;
assign main_genericstandalone_tx_converter_sink_sink_eop = main_genericstandalone_tx_cdc_source_eop;
assign main_genericstandalone_tx_converter_sink_sink_payload_data = main_genericstandalone_tx_cdc_source_payload_data;
assign main_genericstandalone_tx_converter_sink_sink_payload_last_be = main_genericstandalone_tx_cdc_source_payload_last_be;
assign main_genericstandalone_tx_converter_sink_sink_payload_error = main_genericstandalone_tx_cdc_source_payload_error;
assign main_genericstandalone_tx_last_be_sink_stb = main_genericstandalone_tx_converter_source_source_stb;
assign main_genericstandalone_tx_converter_source_source_ack = main_genericstandalone_tx_last_be_sink_ack;
assign main_genericstandalone_tx_last_be_sink_eop = main_genericstandalone_tx_converter_source_source_eop;
assign main_genericstandalone_tx_last_be_sink_payload_data = main_genericstandalone_tx_converter_source_source_payload_data;
assign main_genericstandalone_tx_last_be_sink_payload_last_be = main_genericstandalone_tx_converter_source_source_payload_last_be;
assign main_genericstandalone_tx_last_be_sink_payload_error = main_genericstandalone_tx_converter_source_source_payload_error;
assign main_genericstandalone_padding_inserter_sink_stb = main_genericstandalone_tx_last_be_source_stb;
assign main_genericstandalone_tx_last_be_source_ack = main_genericstandalone_padding_inserter_sink_ack;
assign main_genericstandalone_padding_inserter_sink_eop = main_genericstandalone_tx_last_be_source_eop;
assign main_genericstandalone_padding_inserter_sink_payload_data = main_genericstandalone_tx_last_be_source_payload_data;
assign main_genericstandalone_padding_inserter_sink_payload_last_be = main_genericstandalone_tx_last_be_source_payload_last_be;
assign main_genericstandalone_padding_inserter_sink_payload_error = main_genericstandalone_tx_last_be_source_payload_error;
assign main_genericstandalone_crc32_inserter_sink_stb = main_genericstandalone_padding_inserter_source_stb;
assign main_genericstandalone_padding_inserter_source_ack = main_genericstandalone_crc32_inserter_sink_ack;
assign main_genericstandalone_crc32_inserter_sink_eop = main_genericstandalone_padding_inserter_source_eop;
assign main_genericstandalone_crc32_inserter_sink_payload_data = main_genericstandalone_padding_inserter_source_payload_data;
assign main_genericstandalone_crc32_inserter_sink_payload_last_be = main_genericstandalone_padding_inserter_source_payload_last_be;
assign main_genericstandalone_crc32_inserter_sink_payload_error = main_genericstandalone_padding_inserter_source_payload_error;
assign main_genericstandalone_preamble_inserter_sink_stb = main_genericstandalone_crc32_inserter_source_stb;
assign main_genericstandalone_crc32_inserter_source_ack = main_genericstandalone_preamble_inserter_sink_ack;
assign main_genericstandalone_preamble_inserter_sink_eop = main_genericstandalone_crc32_inserter_source_eop;
assign main_genericstandalone_preamble_inserter_sink_payload_data = main_genericstandalone_crc32_inserter_source_payload_data;
assign main_genericstandalone_preamble_inserter_sink_payload_last_be = main_genericstandalone_crc32_inserter_source_payload_last_be;
assign main_genericstandalone_preamble_inserter_sink_payload_error = main_genericstandalone_crc32_inserter_source_payload_error;
assign main_genericstandalone_tx_gap_inserter_sink_stb = main_genericstandalone_preamble_inserter_source_stb;
assign main_genericstandalone_preamble_inserter_source_ack = main_genericstandalone_tx_gap_inserter_sink_ack;
assign main_genericstandalone_tx_gap_inserter_sink_eop = main_genericstandalone_preamble_inserter_source_eop;
assign main_genericstandalone_tx_gap_inserter_sink_payload_data = main_genericstandalone_preamble_inserter_source_payload_data;
assign main_genericstandalone_tx_gap_inserter_sink_payload_last_be = main_genericstandalone_preamble_inserter_source_payload_last_be;
assign main_genericstandalone_tx_gap_inserter_sink_payload_error = main_genericstandalone_preamble_inserter_source_payload_error;
assign main_genericstandalone_pcs_sink_stb = main_genericstandalone_tx_gap_inserter_source_stb;
assign main_genericstandalone_tx_gap_inserter_source_ack = main_genericstandalone_pcs_sink_ack;
assign main_genericstandalone_pcs_sink_eop = main_genericstandalone_tx_gap_inserter_source_eop;
assign main_genericstandalone_pcs_sink_payload_data = main_genericstandalone_tx_gap_inserter_source_payload_data;
assign main_genericstandalone_pcs_sink_payload_last_be = main_genericstandalone_tx_gap_inserter_source_payload_last_be;
assign main_genericstandalone_pcs_sink_payload_error = main_genericstandalone_tx_gap_inserter_source_payload_error;
assign main_genericstandalone_preamble_checker_sink_stb = main_genericstandalone_pcs_source_stb;
assign main_genericstandalone_pcs_source_ack = main_genericstandalone_preamble_checker_sink_ack;
assign main_genericstandalone_preamble_checker_sink_eop = main_genericstandalone_pcs_source_eop;
assign main_genericstandalone_preamble_checker_sink_payload_data = main_genericstandalone_pcs_source_payload_data;
assign main_genericstandalone_preamble_checker_sink_payload_last_be = main_genericstandalone_pcs_source_payload_last_be;
assign main_genericstandalone_preamble_checker_sink_payload_error = main_genericstandalone_pcs_source_payload_error;
assign main_genericstandalone_crc32_checker_sink_sink_stb = main_genericstandalone_preamble_checker_source_stb;
assign main_genericstandalone_preamble_checker_source_ack = main_genericstandalone_crc32_checker_sink_sink_ack;
assign main_genericstandalone_crc32_checker_sink_sink_eop = main_genericstandalone_preamble_checker_source_eop;
assign main_genericstandalone_crc32_checker_sink_sink_payload_data = main_genericstandalone_preamble_checker_source_payload_data;
assign main_genericstandalone_crc32_checker_sink_sink_payload_last_be = main_genericstandalone_preamble_checker_source_payload_last_be;
assign main_genericstandalone_crc32_checker_sink_sink_payload_error = main_genericstandalone_preamble_checker_source_payload_error;
assign main_genericstandalone_padding_checker_sink_stb = main_genericstandalone_crc32_checker_source_source_stb;
assign main_genericstandalone_crc32_checker_source_source_ack = main_genericstandalone_padding_checker_sink_ack;
assign main_genericstandalone_padding_checker_sink_eop = main_genericstandalone_crc32_checker_source_source_eop;
assign main_genericstandalone_padding_checker_sink_payload_data = main_genericstandalone_crc32_checker_source_source_payload_data;
assign main_genericstandalone_padding_checker_sink_payload_last_be = main_genericstandalone_crc32_checker_source_source_payload_last_be;
assign main_genericstandalone_padding_checker_sink_payload_error = main_genericstandalone_crc32_checker_source_source_payload_error;
assign main_genericstandalone_rx_last_be_sink_stb = main_genericstandalone_padding_checker_source_stb;
assign main_genericstandalone_padding_checker_source_ack = main_genericstandalone_rx_last_be_sink_ack;
assign main_genericstandalone_rx_last_be_sink_eop = main_genericstandalone_padding_checker_source_eop;
assign main_genericstandalone_rx_last_be_sink_payload_data = main_genericstandalone_padding_checker_source_payload_data;
assign main_genericstandalone_rx_last_be_sink_payload_last_be = main_genericstandalone_padding_checker_source_payload_last_be;
assign main_genericstandalone_rx_last_be_sink_payload_error = main_genericstandalone_padding_checker_source_payload_error;
assign main_genericstandalone_rx_converter_sink_sink_stb = main_genericstandalone_rx_last_be_source_stb;
assign main_genericstandalone_rx_last_be_source_ack = main_genericstandalone_rx_converter_sink_sink_ack;
assign main_genericstandalone_rx_converter_sink_sink_eop = main_genericstandalone_rx_last_be_source_eop;
assign main_genericstandalone_rx_converter_sink_sink_payload_data = main_genericstandalone_rx_last_be_source_payload_data;
assign main_genericstandalone_rx_converter_sink_sink_payload_last_be = main_genericstandalone_rx_last_be_source_payload_last_be;
assign main_genericstandalone_rx_converter_sink_sink_payload_error = main_genericstandalone_rx_last_be_source_payload_error;
assign main_genericstandalone_rx_cdc_sink_stb = main_genericstandalone_rx_converter_source_source_stb;
assign main_genericstandalone_rx_converter_source_source_ack = main_genericstandalone_rx_cdc_sink_ack;
assign main_genericstandalone_rx_cdc_sink_eop = main_genericstandalone_rx_converter_source_source_eop;
assign main_genericstandalone_rx_cdc_sink_payload_data = main_genericstandalone_rx_converter_source_source_payload_data;
assign main_genericstandalone_rx_cdc_sink_payload_last_be = main_genericstandalone_rx_converter_source_source_payload_last_be;
assign main_genericstandalone_rx_cdc_sink_payload_error = main_genericstandalone_rx_converter_source_source_payload_error;

// synthesis translate_off
reg dummy_d_35;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_gap_inserter_sink_ack <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_stb <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_eop <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_tx_gap_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_tx_gap_inserter_counter_reset <= 1'd0;
	main_genericstandalone_tx_gap_inserter_counter_ce <= 1'd0;
	builder_liteethmacgap_next_state <= 1'd0;
	builder_liteethmacgap_next_state <= builder_liteethmacgap_state;
	case (builder_liteethmacgap_state)
		1'd1: begin
			main_genericstandalone_tx_gap_inserter_counter_ce <= 1'd1;
			if ((main_genericstandalone_tx_gap_inserter_counter == 4'd11)) begin
				builder_liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_tx_gap_inserter_counter_reset <= 1'd1;
			main_genericstandalone_tx_gap_inserter_source_stb <= main_genericstandalone_tx_gap_inserter_sink_stb;
			main_genericstandalone_tx_gap_inserter_sink_ack <= main_genericstandalone_tx_gap_inserter_source_ack;
			main_genericstandalone_tx_gap_inserter_source_eop <= main_genericstandalone_tx_gap_inserter_sink_eop;
			main_genericstandalone_tx_gap_inserter_source_payload_data <= main_genericstandalone_tx_gap_inserter_sink_payload_data;
			main_genericstandalone_tx_gap_inserter_source_payload_last_be <= main_genericstandalone_tx_gap_inserter_sink_payload_last_be;
			main_genericstandalone_tx_gap_inserter_source_payload_error <= main_genericstandalone_tx_gap_inserter_sink_payload_error;
			if (((main_genericstandalone_tx_gap_inserter_sink_stb & main_genericstandalone_tx_gap_inserter_sink_eop) & main_genericstandalone_tx_gap_inserter_sink_ack)) begin
				builder_liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_35 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_preamble_inserter_source_payload_last_be = main_genericstandalone_preamble_inserter_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_36;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_preamble_inserter_sink_ack <= 1'd0;
	main_genericstandalone_preamble_inserter_source_stb <= 1'd0;
	main_genericstandalone_preamble_inserter_source_eop <= 1'd0;
	main_genericstandalone_preamble_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_preamble_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_preamble_inserter_clr_cnt <= 1'd0;
	main_genericstandalone_preamble_inserter_inc_cnt <= 1'd0;
	builder_liteethmacpreambleinserter_next_state <= 2'd0;
	main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_sink_payload_data;
	builder_liteethmacpreambleinserter_next_state <= builder_liteethmacpreambleinserter_state;
	case (builder_liteethmacpreambleinserter_state)
		1'd1: begin
			main_genericstandalone_preamble_inserter_source_stb <= 1'd1;
			case (main_genericstandalone_preamble_inserter_cnt)
				1'd0: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[55:48];
				end
				default: begin
					main_genericstandalone_preamble_inserter_source_payload_data <= main_genericstandalone_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((main_genericstandalone_preamble_inserter_cnt == 3'd7)) begin
				if (main_genericstandalone_preamble_inserter_source_ack) begin
					builder_liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				main_genericstandalone_preamble_inserter_inc_cnt <= main_genericstandalone_preamble_inserter_source_ack;
			end
		end
		2'd2: begin
			main_genericstandalone_preamble_inserter_source_stb <= main_genericstandalone_preamble_inserter_sink_stb;
			main_genericstandalone_preamble_inserter_sink_ack <= main_genericstandalone_preamble_inserter_source_ack;
			main_genericstandalone_preamble_inserter_source_eop <= main_genericstandalone_preamble_inserter_sink_eop;
			main_genericstandalone_preamble_inserter_source_payload_error <= main_genericstandalone_preamble_inserter_sink_payload_error;
			if (((main_genericstandalone_preamble_inserter_sink_stb & main_genericstandalone_preamble_inserter_sink_eop) & main_genericstandalone_preamble_inserter_source_ack)) begin
				builder_liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_preamble_inserter_sink_ack <= 1'd1;
			main_genericstandalone_preamble_inserter_clr_cnt <= 1'd1;
			if (main_genericstandalone_preamble_inserter_sink_stb) begin
				main_genericstandalone_preamble_inserter_sink_ack <= 1'd0;
				builder_liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_36 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_preamble_checker_source_payload_data = main_genericstandalone_preamble_checker_sink_payload_data;
assign main_genericstandalone_preamble_checker_source_payload_last_be = main_genericstandalone_preamble_checker_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_37;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_preamble_checker_sink_ack <= 1'd0;
	main_genericstandalone_preamble_checker_source_stb <= 1'd0;
	main_genericstandalone_preamble_checker_source_eop <= 1'd0;
	main_genericstandalone_preamble_checker_source_payload_error <= 1'd0;
	main_genericstandalone_preamble_checker_error <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= builder_liteethmacpreamblechecker_state;
	case (builder_liteethmacpreamblechecker_state)
		1'd1: begin
			main_genericstandalone_preamble_checker_source_stb <= main_genericstandalone_preamble_checker_sink_stb;
			main_genericstandalone_preamble_checker_sink_ack <= main_genericstandalone_preamble_checker_source_ack;
			main_genericstandalone_preamble_checker_source_eop <= main_genericstandalone_preamble_checker_sink_eop;
			main_genericstandalone_preamble_checker_source_payload_error <= main_genericstandalone_preamble_checker_sink_payload_error;
			if (((main_genericstandalone_preamble_checker_source_stb & main_genericstandalone_preamble_checker_source_eop) & main_genericstandalone_preamble_checker_source_ack)) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			main_genericstandalone_preamble_checker_sink_ack <= 1'd1;
			if (((main_genericstandalone_preamble_checker_sink_stb & (~main_genericstandalone_preamble_checker_sink_eop)) & (main_genericstandalone_preamble_checker_sink_payload_data == 8'd213))) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((main_genericstandalone_preamble_checker_sink_stb & main_genericstandalone_preamble_checker_sink_eop)) begin
				main_genericstandalone_preamble_checker_error <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_37 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_inserter_cnt_done = (main_genericstandalone_crc32_inserter_cnt == 1'd0);
assign main_genericstandalone_crc32_inserter_data1 = main_genericstandalone_crc32_inserter_data0;
assign main_genericstandalone_crc32_inserter_last = main_genericstandalone_crc32_inserter_reg;
assign main_genericstandalone_crc32_inserter_value = (~{main_genericstandalone_crc32_inserter_reg[0], main_genericstandalone_crc32_inserter_reg[1], main_genericstandalone_crc32_inserter_reg[2], main_genericstandalone_crc32_inserter_reg[3], main_genericstandalone_crc32_inserter_reg[4], main_genericstandalone_crc32_inserter_reg[5], main_genericstandalone_crc32_inserter_reg[6], main_genericstandalone_crc32_inserter_reg[7], main_genericstandalone_crc32_inserter_reg[8], main_genericstandalone_crc32_inserter_reg[9], main_genericstandalone_crc32_inserter_reg[10], main_genericstandalone_crc32_inserter_reg[11], main_genericstandalone_crc32_inserter_reg[12], main_genericstandalone_crc32_inserter_reg[13], main_genericstandalone_crc32_inserter_reg[14], main_genericstandalone_crc32_inserter_reg[15], main_genericstandalone_crc32_inserter_reg[16], main_genericstandalone_crc32_inserter_reg[17], main_genericstandalone_crc32_inserter_reg[18], main_genericstandalone_crc32_inserter_reg[19], main_genericstandalone_crc32_inserter_reg[20], main_genericstandalone_crc32_inserter_reg[21], main_genericstandalone_crc32_inserter_reg[22], main_genericstandalone_crc32_inserter_reg[23], main_genericstandalone_crc32_inserter_reg[24], main_genericstandalone_crc32_inserter_reg[25], main_genericstandalone_crc32_inserter_reg[26], main_genericstandalone_crc32_inserter_reg[27], main_genericstandalone_crc32_inserter_reg[28], main_genericstandalone_crc32_inserter_reg[29], main_genericstandalone_crc32_inserter_reg[30], main_genericstandalone_crc32_inserter_reg[31]});
assign main_genericstandalone_crc32_inserter_error = (main_genericstandalone_crc32_inserter_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_38;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_inserter_next <= 32'd0;
	main_genericstandalone_crc32_inserter_next[0] <= (((main_genericstandalone_crc32_inserter_last[24] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[1] <= (((((((main_genericstandalone_crc32_inserter_last[25] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[2] <= (((((((((main_genericstandalone_crc32_inserter_last[26] ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[3] <= (((((((main_genericstandalone_crc32_inserter_last[27] ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[4] <= (((((((((main_genericstandalone_crc32_inserter_last[28] ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[5] <= (((((((((((((main_genericstandalone_crc32_inserter_last[29] ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[6] <= (((((((((((main_genericstandalone_crc32_inserter_last[30] ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[7] <= (((((((((main_genericstandalone_crc32_inserter_last[31] ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[8] <= ((((((((main_genericstandalone_crc32_inserter_last[0] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[9] <= ((((((((main_genericstandalone_crc32_inserter_last[1] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[10] <= ((((((((main_genericstandalone_crc32_inserter_last[2] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[11] <= ((((((((main_genericstandalone_crc32_inserter_last[3] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[12] <= ((((((((((((main_genericstandalone_crc32_inserter_last[4] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[13] <= ((((((((((((main_genericstandalone_crc32_inserter_last[5] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[14] <= ((((((((((main_genericstandalone_crc32_inserter_last[6] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[15] <= ((((((((main_genericstandalone_crc32_inserter_last[7] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[16] <= ((((((main_genericstandalone_crc32_inserter_last[8] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[17] <= ((((((main_genericstandalone_crc32_inserter_last[9] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[18] <= ((((((main_genericstandalone_crc32_inserter_last[10] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[19] <= ((((main_genericstandalone_crc32_inserter_last[11] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[20] <= ((main_genericstandalone_crc32_inserter_last[12] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]);
	main_genericstandalone_crc32_inserter_next[21] <= ((main_genericstandalone_crc32_inserter_last[13] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]);
	main_genericstandalone_crc32_inserter_next[22] <= ((main_genericstandalone_crc32_inserter_last[14] ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[23] <= ((((((main_genericstandalone_crc32_inserter_last[15] ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_data1[6]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[24] <= ((((((main_genericstandalone_crc32_inserter_last[16] ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[25] <= ((((main_genericstandalone_crc32_inserter_last[17] ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[26] <= ((((((((main_genericstandalone_crc32_inserter_last[18] ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]) ^ main_genericstandalone_crc32_inserter_last[24]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_data1[7]);
	main_genericstandalone_crc32_inserter_next[27] <= ((((((((main_genericstandalone_crc32_inserter_last[19] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]) ^ main_genericstandalone_crc32_inserter_last[25]) ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_data1[6]);
	main_genericstandalone_crc32_inserter_next[28] <= ((((((main_genericstandalone_crc32_inserter_last[20] ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]) ^ main_genericstandalone_crc32_inserter_last[26]) ^ main_genericstandalone_crc32_inserter_data1[5]);
	main_genericstandalone_crc32_inserter_next[29] <= ((((((main_genericstandalone_crc32_inserter_last[21] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[30]) ^ main_genericstandalone_crc32_inserter_data1[1]) ^ main_genericstandalone_crc32_inserter_last[27]) ^ main_genericstandalone_crc32_inserter_data1[4]);
	main_genericstandalone_crc32_inserter_next[30] <= ((((main_genericstandalone_crc32_inserter_last[22] ^ main_genericstandalone_crc32_inserter_last[31]) ^ main_genericstandalone_crc32_inserter_data1[0]) ^ main_genericstandalone_crc32_inserter_last[28]) ^ main_genericstandalone_crc32_inserter_data1[3]);
	main_genericstandalone_crc32_inserter_next[31] <= ((main_genericstandalone_crc32_inserter_last[23] ^ main_genericstandalone_crc32_inserter_last[29]) ^ main_genericstandalone_crc32_inserter_data1[2]);
// synthesis translate_off
	dummy_d_38 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_39;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_inserter_sink_ack <= 1'd0;
	main_genericstandalone_crc32_inserter_source_stb <= 1'd0;
	main_genericstandalone_crc32_inserter_source_eop <= 1'd0;
	main_genericstandalone_crc32_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_crc32_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_crc32_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_crc32_inserter_data0 <= 8'd0;
	main_genericstandalone_crc32_inserter_ce <= 1'd0;
	main_genericstandalone_crc32_inserter_reset <= 1'd0;
	main_genericstandalone_crc32_inserter_is_ongoing0 <= 1'd0;
	main_genericstandalone_crc32_inserter_is_ongoing1 <= 1'd0;
	builder_liteethmaccrc32inserter_next_state <= 2'd0;
	builder_liteethmaccrc32inserter_next_state <= builder_liteethmaccrc32inserter_state;
	case (builder_liteethmaccrc32inserter_state)
		1'd1: begin
			main_genericstandalone_crc32_inserter_ce <= (main_genericstandalone_crc32_inserter_sink_stb & main_genericstandalone_crc32_inserter_source_ack);
			main_genericstandalone_crc32_inserter_data0 <= main_genericstandalone_crc32_inserter_sink_payload_data;
			main_genericstandalone_crc32_inserter_source_stb <= main_genericstandalone_crc32_inserter_sink_stb;
			main_genericstandalone_crc32_inserter_sink_ack <= main_genericstandalone_crc32_inserter_source_ack;
			main_genericstandalone_crc32_inserter_source_eop <= main_genericstandalone_crc32_inserter_sink_eop;
			main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_sink_payload_data;
			main_genericstandalone_crc32_inserter_source_payload_last_be <= main_genericstandalone_crc32_inserter_sink_payload_last_be;
			main_genericstandalone_crc32_inserter_source_payload_error <= main_genericstandalone_crc32_inserter_sink_payload_error;
			main_genericstandalone_crc32_inserter_source_eop <= 1'd0;
			if (((main_genericstandalone_crc32_inserter_sink_stb & main_genericstandalone_crc32_inserter_sink_eop) & main_genericstandalone_crc32_inserter_source_ack)) begin
				builder_liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_genericstandalone_crc32_inserter_source_stb <= 1'd1;
			case (main_genericstandalone_crc32_inserter_cnt)
				1'd0: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[31:24];
				end
				1'd1: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[23:16];
				end
				2'd2: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[15:8];
				end
				default: begin
					main_genericstandalone_crc32_inserter_source_payload_data <= main_genericstandalone_crc32_inserter_value[7:0];
				end
			endcase
			if (main_genericstandalone_crc32_inserter_cnt_done) begin
				main_genericstandalone_crc32_inserter_source_eop <= 1'd1;
				if (main_genericstandalone_crc32_inserter_source_ack) begin
					builder_liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			main_genericstandalone_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			main_genericstandalone_crc32_inserter_reset <= 1'd1;
			main_genericstandalone_crc32_inserter_sink_ack <= 1'd1;
			if (main_genericstandalone_crc32_inserter_sink_stb) begin
				main_genericstandalone_crc32_inserter_sink_ack <= 1'd0;
				builder_liteethmaccrc32inserter_next_state <= 1'd1;
			end
			main_genericstandalone_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_39 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_fifo_full = (main_genericstandalone_crc32_checker_syncfifo_level == 3'd4);
assign main_genericstandalone_crc32_checker_fifo_in = (main_genericstandalone_crc32_checker_sink_sink_stb & ((~main_genericstandalone_crc32_checker_fifo_full) | main_genericstandalone_crc32_checker_fifo_out));
assign main_genericstandalone_crc32_checker_fifo_out = (main_genericstandalone_crc32_checker_source_source_stb & main_genericstandalone_crc32_checker_source_source_ack);
assign main_genericstandalone_crc32_checker_syncfifo_sink_eop = main_genericstandalone_crc32_checker_sink_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_data = main_genericstandalone_crc32_checker_sink_sink_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be = main_genericstandalone_crc32_checker_sink_sink_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_sink_payload_error = main_genericstandalone_crc32_checker_sink_sink_payload_error;

// synthesis translate_off
reg dummy_d_40;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= 1'd0;
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= main_genericstandalone_crc32_checker_sink_sink_stb;
	main_genericstandalone_crc32_checker_syncfifo_sink_stb <= main_genericstandalone_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_40 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_41;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_sink_sink_ack <= 1'd0;
	main_genericstandalone_crc32_checker_sink_sink_ack <= main_genericstandalone_crc32_checker_syncfifo_sink_ack;
	main_genericstandalone_crc32_checker_sink_sink_ack <= main_genericstandalone_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_41 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_source_source_stb = (main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_fifo_full);
assign main_genericstandalone_crc32_checker_source_source_eop = main_genericstandalone_crc32_checker_sink_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_source_ack = main_genericstandalone_crc32_checker_fifo_out;
assign main_genericstandalone_crc32_checker_source_source_payload_data = main_genericstandalone_crc32_checker_syncfifo_source_payload_data;
assign main_genericstandalone_crc32_checker_source_source_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be;

// synthesis translate_off
reg dummy_d_42;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_source_source_payload_error <= 1'd0;
	main_genericstandalone_crc32_checker_source_source_payload_error <= main_genericstandalone_crc32_checker_syncfifo_source_payload_error;
	main_genericstandalone_crc32_checker_source_source_payload_error <= (main_genericstandalone_crc32_checker_sink_sink_payload_error | main_genericstandalone_crc32_checker_crc_error);
// synthesis translate_off
	dummy_d_42 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_error = ((main_genericstandalone_crc32_checker_source_source_stb & main_genericstandalone_crc32_checker_source_source_eop) & main_genericstandalone_crc32_checker_crc_error);
assign main_genericstandalone_crc32_checker_crc_data0 = main_genericstandalone_crc32_checker_sink_sink_payload_data;
assign main_genericstandalone_crc32_checker_crc_data1 = main_genericstandalone_crc32_checker_crc_data0;
assign main_genericstandalone_crc32_checker_crc_last = main_genericstandalone_crc32_checker_crc_reg;
assign main_genericstandalone_crc32_checker_crc_value = (~{main_genericstandalone_crc32_checker_crc_reg[0], main_genericstandalone_crc32_checker_crc_reg[1], main_genericstandalone_crc32_checker_crc_reg[2], main_genericstandalone_crc32_checker_crc_reg[3], main_genericstandalone_crc32_checker_crc_reg[4], main_genericstandalone_crc32_checker_crc_reg[5], main_genericstandalone_crc32_checker_crc_reg[6], main_genericstandalone_crc32_checker_crc_reg[7], main_genericstandalone_crc32_checker_crc_reg[8], main_genericstandalone_crc32_checker_crc_reg[9], main_genericstandalone_crc32_checker_crc_reg[10], main_genericstandalone_crc32_checker_crc_reg[11], main_genericstandalone_crc32_checker_crc_reg[12], main_genericstandalone_crc32_checker_crc_reg[13], main_genericstandalone_crc32_checker_crc_reg[14], main_genericstandalone_crc32_checker_crc_reg[15], main_genericstandalone_crc32_checker_crc_reg[16], main_genericstandalone_crc32_checker_crc_reg[17], main_genericstandalone_crc32_checker_crc_reg[18], main_genericstandalone_crc32_checker_crc_reg[19], main_genericstandalone_crc32_checker_crc_reg[20], main_genericstandalone_crc32_checker_crc_reg[21], main_genericstandalone_crc32_checker_crc_reg[22], main_genericstandalone_crc32_checker_crc_reg[23], main_genericstandalone_crc32_checker_crc_reg[24], main_genericstandalone_crc32_checker_crc_reg[25], main_genericstandalone_crc32_checker_crc_reg[26], main_genericstandalone_crc32_checker_crc_reg[27], main_genericstandalone_crc32_checker_crc_reg[28], main_genericstandalone_crc32_checker_crc_reg[29], main_genericstandalone_crc32_checker_crc_reg[30], main_genericstandalone_crc32_checker_crc_reg[31]});
assign main_genericstandalone_crc32_checker_crc_error = (main_genericstandalone_crc32_checker_crc_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_43;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_crc_next <= 32'd0;
	main_genericstandalone_crc32_checker_crc_next[0] <= (((main_genericstandalone_crc32_checker_crc_last[24] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[1] <= (((((((main_genericstandalone_crc32_checker_crc_last[25] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[2] <= (((((((((main_genericstandalone_crc32_checker_crc_last[26] ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[3] <= (((((((main_genericstandalone_crc32_checker_crc_last[27] ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[4] <= (((((((((main_genericstandalone_crc32_checker_crc_last[28] ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[5] <= (((((((((((((main_genericstandalone_crc32_checker_crc_last[29] ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[6] <= (((((((((((main_genericstandalone_crc32_checker_crc_last[30] ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[7] <= (((((((((main_genericstandalone_crc32_checker_crc_last[31] ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[8] <= ((((((((main_genericstandalone_crc32_checker_crc_last[0] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[9] <= ((((((((main_genericstandalone_crc32_checker_crc_last[1] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[10] <= ((((((((main_genericstandalone_crc32_checker_crc_last[2] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[11] <= ((((((((main_genericstandalone_crc32_checker_crc_last[3] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[12] <= ((((((((((((main_genericstandalone_crc32_checker_crc_last[4] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[13] <= ((((((((((((main_genericstandalone_crc32_checker_crc_last[5] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[14] <= ((((((((((main_genericstandalone_crc32_checker_crc_last[6] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[15] <= ((((((((main_genericstandalone_crc32_checker_crc_last[7] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[16] <= ((((((main_genericstandalone_crc32_checker_crc_last[8] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[17] <= ((((((main_genericstandalone_crc32_checker_crc_last[9] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[18] <= ((((((main_genericstandalone_crc32_checker_crc_last[10] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[19] <= ((((main_genericstandalone_crc32_checker_crc_last[11] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[20] <= ((main_genericstandalone_crc32_checker_crc_last[12] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]);
	main_genericstandalone_crc32_checker_crc_next[21] <= ((main_genericstandalone_crc32_checker_crc_last[13] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]);
	main_genericstandalone_crc32_checker_crc_next[22] <= ((main_genericstandalone_crc32_checker_crc_last[14] ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[23] <= ((((((main_genericstandalone_crc32_checker_crc_last[15] ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_data1[6]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[24] <= ((((((main_genericstandalone_crc32_checker_crc_last[16] ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[25] <= ((((main_genericstandalone_crc32_checker_crc_last[17] ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[26] <= ((((((((main_genericstandalone_crc32_checker_crc_last[18] ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]) ^ main_genericstandalone_crc32_checker_crc_last[24]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_data1[7]);
	main_genericstandalone_crc32_checker_crc_next[27] <= ((((((((main_genericstandalone_crc32_checker_crc_last[19] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]) ^ main_genericstandalone_crc32_checker_crc_last[25]) ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_data1[6]);
	main_genericstandalone_crc32_checker_crc_next[28] <= ((((((main_genericstandalone_crc32_checker_crc_last[20] ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]) ^ main_genericstandalone_crc32_checker_crc_last[26]) ^ main_genericstandalone_crc32_checker_crc_data1[5]);
	main_genericstandalone_crc32_checker_crc_next[29] <= ((((((main_genericstandalone_crc32_checker_crc_last[21] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[30]) ^ main_genericstandalone_crc32_checker_crc_data1[1]) ^ main_genericstandalone_crc32_checker_crc_last[27]) ^ main_genericstandalone_crc32_checker_crc_data1[4]);
	main_genericstandalone_crc32_checker_crc_next[30] <= ((((main_genericstandalone_crc32_checker_crc_last[22] ^ main_genericstandalone_crc32_checker_crc_last[31]) ^ main_genericstandalone_crc32_checker_crc_data1[0]) ^ main_genericstandalone_crc32_checker_crc_last[28]) ^ main_genericstandalone_crc32_checker_crc_data1[3]);
	main_genericstandalone_crc32_checker_crc_next[31] <= ((main_genericstandalone_crc32_checker_crc_last[23] ^ main_genericstandalone_crc32_checker_crc_last[29]) ^ main_genericstandalone_crc32_checker_crc_data1[2]);
// synthesis translate_off
	dummy_d_43 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_din = {main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be, main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data};
assign {main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be, main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data} = main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout;
assign main_genericstandalone_crc32_checker_syncfifo_sink_ack = main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_we = main_genericstandalone_crc32_checker_syncfifo_sink_stb;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_eop = main_genericstandalone_crc32_checker_syncfifo_sink_eop;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_data = main_genericstandalone_crc32_checker_syncfifo_sink_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_sink_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_fifo_in_payload_error = main_genericstandalone_crc32_checker_syncfifo_sink_payload_error;
assign main_genericstandalone_crc32_checker_syncfifo_source_stb = main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable;
assign main_genericstandalone_crc32_checker_syncfifo_source_eop = main_genericstandalone_crc32_checker_syncfifo_fifo_out_eop;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_data = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_data;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_last_be = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign main_genericstandalone_crc32_checker_syncfifo_source_payload_error = main_genericstandalone_crc32_checker_syncfifo_fifo_out_payload_error;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_re = main_genericstandalone_crc32_checker_syncfifo_source_ack;

// synthesis translate_off
reg dummy_d_44;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (main_genericstandalone_crc32_checker_syncfifo_replace) begin
		main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= (main_genericstandalone_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		main_genericstandalone_crc32_checker_syncfifo_wrport_adr <= main_genericstandalone_crc32_checker_syncfifo_produce;
	end
// synthesis translate_off
	dummy_d_44 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w = main_genericstandalone_crc32_checker_syncfifo_syncfifo_din;
assign main_genericstandalone_crc32_checker_syncfifo_wrport_we = (main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & (main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable | main_genericstandalone_crc32_checker_syncfifo_replace));
assign main_genericstandalone_crc32_checker_syncfifo_do_read = (main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable & main_genericstandalone_crc32_checker_syncfifo_syncfifo_re);
assign main_genericstandalone_crc32_checker_syncfifo_rdport_adr = main_genericstandalone_crc32_checker_syncfifo_consume;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_dout = main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r;
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable = (main_genericstandalone_crc32_checker_syncfifo_level != 3'd5);
assign main_genericstandalone_crc32_checker_syncfifo_syncfifo_readable = (main_genericstandalone_crc32_checker_syncfifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_45;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_crc32_checker_crc_ce <= 1'd0;
	main_genericstandalone_crc32_checker_crc_reset <= 1'd0;
	main_genericstandalone_crc32_checker_fifo_reset <= 1'd0;
	builder_liteethmaccrc32checker_next_state <= 2'd0;
	builder_liteethmaccrc32checker_next_state <= builder_liteethmaccrc32checker_state;
	case (builder_liteethmaccrc32checker_state)
		1'd1: begin
			if ((main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_sink_sink_ack)) begin
				main_genericstandalone_crc32_checker_crc_ce <= 1'd1;
				builder_liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((main_genericstandalone_crc32_checker_sink_sink_stb & main_genericstandalone_crc32_checker_sink_sink_ack)) begin
				main_genericstandalone_crc32_checker_crc_ce <= 1'd1;
				if (main_genericstandalone_crc32_checker_sink_sink_eop) begin
					builder_liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_genericstandalone_crc32_checker_crc_reset <= 1'd1;
			main_genericstandalone_crc32_checker_fifo_reset <= 1'd1;
			builder_liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_45 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_ps_preamble_error_o = (main_genericstandalone_ps_preamble_error_toggle_o ^ main_genericstandalone_ps_preamble_error_toggle_o_r);
assign main_genericstandalone_ps_crc_error_o = (main_genericstandalone_ps_crc_error_toggle_o ^ main_genericstandalone_ps_crc_error_toggle_o_r);
assign main_genericstandalone_padding_inserter_counter_done = (main_genericstandalone_padding_inserter_counter >= 6'd59);

// synthesis translate_off
reg dummy_d_46;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_padding_inserter_sink_ack <= 1'd0;
	main_genericstandalone_padding_inserter_source_stb <= 1'd0;
	main_genericstandalone_padding_inserter_source_eop <= 1'd0;
	main_genericstandalone_padding_inserter_source_payload_data <= 8'd0;
	main_genericstandalone_padding_inserter_source_payload_last_be <= 1'd0;
	main_genericstandalone_padding_inserter_source_payload_error <= 1'd0;
	main_genericstandalone_padding_inserter_counter_reset <= 1'd0;
	main_genericstandalone_padding_inserter_counter_ce <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= builder_liteethmacpaddinginserter_state;
	case (builder_liteethmacpaddinginserter_state)
		1'd1: begin
			main_genericstandalone_padding_inserter_source_stb <= 1'd1;
			main_genericstandalone_padding_inserter_source_eop <= main_genericstandalone_padding_inserter_counter_done;
			main_genericstandalone_padding_inserter_source_payload_data <= 1'd0;
			if ((main_genericstandalone_padding_inserter_source_stb & main_genericstandalone_padding_inserter_source_ack)) begin
				main_genericstandalone_padding_inserter_counter_ce <= 1'd1;
				if (main_genericstandalone_padding_inserter_counter_done) begin
					main_genericstandalone_padding_inserter_counter_reset <= 1'd1;
					builder_liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_genericstandalone_padding_inserter_source_stb <= main_genericstandalone_padding_inserter_sink_stb;
			main_genericstandalone_padding_inserter_sink_ack <= main_genericstandalone_padding_inserter_source_ack;
			main_genericstandalone_padding_inserter_source_eop <= main_genericstandalone_padding_inserter_sink_eop;
			main_genericstandalone_padding_inserter_source_payload_data <= main_genericstandalone_padding_inserter_sink_payload_data;
			main_genericstandalone_padding_inserter_source_payload_last_be <= main_genericstandalone_padding_inserter_sink_payload_last_be;
			main_genericstandalone_padding_inserter_source_payload_error <= main_genericstandalone_padding_inserter_sink_payload_error;
			if ((main_genericstandalone_padding_inserter_source_stb & main_genericstandalone_padding_inserter_source_ack)) begin
				main_genericstandalone_padding_inserter_counter_ce <= 1'd1;
				if (main_genericstandalone_padding_inserter_sink_eop) begin
					if ((~main_genericstandalone_padding_inserter_counter_done)) begin
						main_genericstandalone_padding_inserter_source_eop <= 1'd0;
						builder_liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						main_genericstandalone_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_46 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_padding_checker_source_stb = main_genericstandalone_padding_checker_sink_stb;
assign main_genericstandalone_padding_checker_sink_ack = main_genericstandalone_padding_checker_source_ack;
assign main_genericstandalone_padding_checker_source_eop = main_genericstandalone_padding_checker_sink_eop;
assign main_genericstandalone_padding_checker_source_payload_data = main_genericstandalone_padding_checker_sink_payload_data;
assign main_genericstandalone_padding_checker_source_payload_last_be = main_genericstandalone_padding_checker_sink_payload_last_be;
assign main_genericstandalone_padding_checker_source_payload_error = main_genericstandalone_padding_checker_sink_payload_error;
assign main_genericstandalone_tx_last_be_source_stb = (main_genericstandalone_tx_last_be_sink_stb & main_genericstandalone_tx_last_be_ongoing);
assign main_genericstandalone_tx_last_be_source_eop = main_genericstandalone_tx_last_be_sink_payload_last_be;
assign main_genericstandalone_tx_last_be_source_payload_data = main_genericstandalone_tx_last_be_sink_payload_data;
assign main_genericstandalone_tx_last_be_sink_ack = main_genericstandalone_tx_last_be_source_ack;
assign main_genericstandalone_rx_last_be_source_stb = main_genericstandalone_rx_last_be_sink_stb;
assign main_genericstandalone_rx_last_be_sink_ack = main_genericstandalone_rx_last_be_source_ack;
assign main_genericstandalone_rx_last_be_source_eop = main_genericstandalone_rx_last_be_sink_eop;
assign main_genericstandalone_rx_last_be_source_payload_data = main_genericstandalone_rx_last_be_sink_payload_data;
assign main_genericstandalone_rx_last_be_source_payload_error = main_genericstandalone_rx_last_be_sink_payload_error;

// synthesis translate_off
reg dummy_d_47;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_last_be_source_payload_last_be <= 1'd0;
	main_genericstandalone_rx_last_be_source_payload_last_be <= main_genericstandalone_rx_last_be_sink_payload_last_be;
	main_genericstandalone_rx_last_be_source_payload_last_be <= main_genericstandalone_rx_last_be_sink_eop;
// synthesis translate_off
	dummy_d_47 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_converter_converter_sink_stb = main_genericstandalone_tx_converter_sink_sink_stb;
assign main_genericstandalone_tx_converter_converter_sink_eop = main_genericstandalone_tx_converter_sink_sink_eop;
assign main_genericstandalone_tx_converter_sink_sink_ack = main_genericstandalone_tx_converter_converter_sink_ack;

// synthesis translate_off
reg dummy_d_48;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_converter_converter_sink_payload_data <= 40'd0;
	main_genericstandalone_tx_converter_converter_sink_payload_data[7:0] <= main_genericstandalone_tx_converter_sink_sink_payload_data[7:0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[8] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[9] <= main_genericstandalone_tx_converter_sink_sink_payload_error[0];
	main_genericstandalone_tx_converter_converter_sink_payload_data[17:10] <= main_genericstandalone_tx_converter_sink_sink_payload_data[15:8];
	main_genericstandalone_tx_converter_converter_sink_payload_data[18] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[1];
	main_genericstandalone_tx_converter_converter_sink_payload_data[19] <= main_genericstandalone_tx_converter_sink_sink_payload_error[1];
	main_genericstandalone_tx_converter_converter_sink_payload_data[27:20] <= main_genericstandalone_tx_converter_sink_sink_payload_data[23:16];
	main_genericstandalone_tx_converter_converter_sink_payload_data[28] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[2];
	main_genericstandalone_tx_converter_converter_sink_payload_data[29] <= main_genericstandalone_tx_converter_sink_sink_payload_error[2];
	main_genericstandalone_tx_converter_converter_sink_payload_data[37:30] <= main_genericstandalone_tx_converter_sink_sink_payload_data[31:24];
	main_genericstandalone_tx_converter_converter_sink_payload_data[38] <= main_genericstandalone_tx_converter_sink_sink_payload_last_be[3];
	main_genericstandalone_tx_converter_converter_sink_payload_data[39] <= main_genericstandalone_tx_converter_sink_sink_payload_error[3];
// synthesis translate_off
	dummy_d_48 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_converter_source_source_stb = main_genericstandalone_tx_converter_converter_source_stb;
assign main_genericstandalone_tx_converter_source_source_eop = main_genericstandalone_tx_converter_converter_source_eop;
assign main_genericstandalone_tx_converter_converter_source_ack = main_genericstandalone_tx_converter_source_source_ack;
assign {main_genericstandalone_tx_converter_source_source_payload_error, main_genericstandalone_tx_converter_source_source_payload_last_be, main_genericstandalone_tx_converter_source_source_payload_data} = main_genericstandalone_tx_converter_converter_source_payload_data;
assign main_genericstandalone_tx_converter_converter_last = (main_genericstandalone_tx_converter_converter_mux == 2'd3);
assign main_genericstandalone_tx_converter_converter_source_stb = main_genericstandalone_tx_converter_converter_sink_stb;
assign main_genericstandalone_tx_converter_converter_source_eop = (main_genericstandalone_tx_converter_converter_sink_eop & main_genericstandalone_tx_converter_converter_last);
assign main_genericstandalone_tx_converter_converter_sink_ack = (main_genericstandalone_tx_converter_converter_last & main_genericstandalone_tx_converter_converter_source_ack);

// synthesis translate_off
reg dummy_d_49;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_converter_converter_source_payload_data <= 10'd0;
	case (main_genericstandalone_tx_converter_converter_mux)
		1'd0: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[39:30];
		end
		1'd1: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd2: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[19:10];
		end
		default: begin
			main_genericstandalone_tx_converter_converter_source_payload_data <= main_genericstandalone_tx_converter_converter_sink_payload_data[9:0];
		end
	endcase
// synthesis translate_off
	dummy_d_49 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_converter_converter_sink_stb = main_genericstandalone_rx_converter_sink_sink_stb;
assign main_genericstandalone_rx_converter_converter_sink_eop = main_genericstandalone_rx_converter_sink_sink_eop;
assign main_genericstandalone_rx_converter_sink_sink_ack = main_genericstandalone_rx_converter_converter_sink_ack;
assign main_genericstandalone_rx_converter_converter_sink_payload_data = {main_genericstandalone_rx_converter_sink_sink_payload_error, main_genericstandalone_rx_converter_sink_sink_payload_last_be, main_genericstandalone_rx_converter_sink_sink_payload_data};
assign main_genericstandalone_rx_converter_source_source_stb = main_genericstandalone_rx_converter_converter_source_stb;
assign main_genericstandalone_rx_converter_source_source_eop = main_genericstandalone_rx_converter_converter_source_eop;
assign main_genericstandalone_rx_converter_converter_source_ack = main_genericstandalone_rx_converter_source_source_ack;

// synthesis translate_off
reg dummy_d_50;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_data <= 32'd0;
	main_genericstandalone_rx_converter_source_source_payload_data[7:0] <= main_genericstandalone_rx_converter_converter_source_payload_data[7:0];
	main_genericstandalone_rx_converter_source_source_payload_data[15:8] <= main_genericstandalone_rx_converter_converter_source_payload_data[17:10];
	main_genericstandalone_rx_converter_source_source_payload_data[23:16] <= main_genericstandalone_rx_converter_converter_source_payload_data[27:20];
	main_genericstandalone_rx_converter_source_source_payload_data[31:24] <= main_genericstandalone_rx_converter_converter_source_payload_data[37:30];
// synthesis translate_off
	dummy_d_50 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_51;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_last_be <= 4'd0;
	main_genericstandalone_rx_converter_source_source_payload_last_be[0] <= main_genericstandalone_rx_converter_converter_source_payload_data[8];
	main_genericstandalone_rx_converter_source_source_payload_last_be[1] <= main_genericstandalone_rx_converter_converter_source_payload_data[18];
	main_genericstandalone_rx_converter_source_source_payload_last_be[2] <= main_genericstandalone_rx_converter_converter_source_payload_data[28];
	main_genericstandalone_rx_converter_source_source_payload_last_be[3] <= main_genericstandalone_rx_converter_converter_source_payload_data[38];
// synthesis translate_off
	dummy_d_51 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_52;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_converter_source_source_payload_error <= 4'd0;
	main_genericstandalone_rx_converter_source_source_payload_error[0] <= main_genericstandalone_rx_converter_converter_source_payload_data[9];
	main_genericstandalone_rx_converter_source_source_payload_error[1] <= main_genericstandalone_rx_converter_converter_source_payload_data[19];
	main_genericstandalone_rx_converter_source_source_payload_error[2] <= main_genericstandalone_rx_converter_converter_source_payload_data[29];
	main_genericstandalone_rx_converter_source_source_payload_error[3] <= main_genericstandalone_rx_converter_converter_source_payload_data[39];
// synthesis translate_off
	dummy_d_52 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_converter_converter_sink_ack = ((~main_genericstandalone_rx_converter_converter_strobe_all) | main_genericstandalone_rx_converter_converter_source_ack);
assign main_genericstandalone_rx_converter_converter_source_stb = main_genericstandalone_rx_converter_converter_strobe_all;
assign main_genericstandalone_rx_converter_converter_load_part = (main_genericstandalone_rx_converter_converter_sink_stb & main_genericstandalone_rx_converter_converter_sink_ack);
assign main_genericstandalone_tx_cdc_asyncfifo_din = {main_genericstandalone_tx_cdc_fifo_in_eop, main_genericstandalone_tx_cdc_fifo_in_payload_error, main_genericstandalone_tx_cdc_fifo_in_payload_last_be, main_genericstandalone_tx_cdc_fifo_in_payload_data};
assign {main_genericstandalone_tx_cdc_fifo_out_eop, main_genericstandalone_tx_cdc_fifo_out_payload_error, main_genericstandalone_tx_cdc_fifo_out_payload_last_be, main_genericstandalone_tx_cdc_fifo_out_payload_data} = main_genericstandalone_tx_cdc_asyncfifo_dout;
assign main_genericstandalone_tx_cdc_sink_ack = main_genericstandalone_tx_cdc_asyncfifo_writable;
assign main_genericstandalone_tx_cdc_asyncfifo_we = main_genericstandalone_tx_cdc_sink_stb;
assign main_genericstandalone_tx_cdc_fifo_in_eop = main_genericstandalone_tx_cdc_sink_eop;
assign main_genericstandalone_tx_cdc_fifo_in_payload_data = main_genericstandalone_tx_cdc_sink_payload_data;
assign main_genericstandalone_tx_cdc_fifo_in_payload_last_be = main_genericstandalone_tx_cdc_sink_payload_last_be;
assign main_genericstandalone_tx_cdc_fifo_in_payload_error = main_genericstandalone_tx_cdc_sink_payload_error;
assign main_genericstandalone_tx_cdc_source_stb = main_genericstandalone_tx_cdc_asyncfifo_readable;
assign main_genericstandalone_tx_cdc_source_eop = main_genericstandalone_tx_cdc_fifo_out_eop;
assign main_genericstandalone_tx_cdc_source_payload_data = main_genericstandalone_tx_cdc_fifo_out_payload_data;
assign main_genericstandalone_tx_cdc_source_payload_last_be = main_genericstandalone_tx_cdc_fifo_out_payload_last_be;
assign main_genericstandalone_tx_cdc_source_payload_error = main_genericstandalone_tx_cdc_fifo_out_payload_error;
assign main_genericstandalone_tx_cdc_asyncfifo_re = main_genericstandalone_tx_cdc_source_ack;
assign main_genericstandalone_tx_cdc_graycounter0_ce = (main_genericstandalone_tx_cdc_asyncfifo_writable & main_genericstandalone_tx_cdc_asyncfifo_we);
assign main_genericstandalone_tx_cdc_graycounter1_ce = (main_genericstandalone_tx_cdc_asyncfifo_readable & main_genericstandalone_tx_cdc_asyncfifo_re);
assign main_genericstandalone_tx_cdc_asyncfifo_writable = (((main_genericstandalone_tx_cdc_graycounter0_q[6] == main_genericstandalone_tx_cdc_consume_wdomain[6]) | (main_genericstandalone_tx_cdc_graycounter0_q[5] == main_genericstandalone_tx_cdc_consume_wdomain[5])) | (main_genericstandalone_tx_cdc_graycounter0_q[4:0] != main_genericstandalone_tx_cdc_consume_wdomain[4:0]));
assign main_genericstandalone_tx_cdc_asyncfifo_readable = (main_genericstandalone_tx_cdc_graycounter1_q != main_genericstandalone_tx_cdc_produce_rdomain);
assign main_genericstandalone_tx_cdc_wrport_adr = main_genericstandalone_tx_cdc_graycounter0_q_binary[5:0];
assign main_genericstandalone_tx_cdc_wrport_dat_w = main_genericstandalone_tx_cdc_asyncfifo_din;
assign main_genericstandalone_tx_cdc_wrport_we = main_genericstandalone_tx_cdc_graycounter0_ce;
assign main_genericstandalone_tx_cdc_rdport_adr = main_genericstandalone_tx_cdc_graycounter1_q_next_binary[5:0];
assign main_genericstandalone_tx_cdc_asyncfifo_dout = main_genericstandalone_tx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_53;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_genericstandalone_tx_cdc_graycounter0_ce) begin
		main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= (main_genericstandalone_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_genericstandalone_tx_cdc_graycounter0_q_next_binary <= main_genericstandalone_tx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_53 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_cdc_graycounter0_q_next = (main_genericstandalone_tx_cdc_graycounter0_q_next_binary ^ main_genericstandalone_tx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_54;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_genericstandalone_tx_cdc_graycounter1_ce) begin
		main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= (main_genericstandalone_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_genericstandalone_tx_cdc_graycounter1_q_next_binary <= main_genericstandalone_tx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_54 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_tx_cdc_graycounter1_q_next = (main_genericstandalone_tx_cdc_graycounter1_q_next_binary ^ main_genericstandalone_tx_cdc_graycounter1_q_next_binary[6:1]);
assign main_genericstandalone_rx_cdc_asyncfifo_din = {main_genericstandalone_rx_cdc_fifo_in_eop, main_genericstandalone_rx_cdc_fifo_in_payload_error, main_genericstandalone_rx_cdc_fifo_in_payload_last_be, main_genericstandalone_rx_cdc_fifo_in_payload_data};
assign {main_genericstandalone_rx_cdc_fifo_out_eop, main_genericstandalone_rx_cdc_fifo_out_payload_error, main_genericstandalone_rx_cdc_fifo_out_payload_last_be, main_genericstandalone_rx_cdc_fifo_out_payload_data} = main_genericstandalone_rx_cdc_asyncfifo_dout;
assign main_genericstandalone_rx_cdc_sink_ack = main_genericstandalone_rx_cdc_asyncfifo_writable;
assign main_genericstandalone_rx_cdc_asyncfifo_we = main_genericstandalone_rx_cdc_sink_stb;
assign main_genericstandalone_rx_cdc_fifo_in_eop = main_genericstandalone_rx_cdc_sink_eop;
assign main_genericstandalone_rx_cdc_fifo_in_payload_data = main_genericstandalone_rx_cdc_sink_payload_data;
assign main_genericstandalone_rx_cdc_fifo_in_payload_last_be = main_genericstandalone_rx_cdc_sink_payload_last_be;
assign main_genericstandalone_rx_cdc_fifo_in_payload_error = main_genericstandalone_rx_cdc_sink_payload_error;
assign main_genericstandalone_rx_cdc_source_stb = main_genericstandalone_rx_cdc_asyncfifo_readable;
assign main_genericstandalone_rx_cdc_source_eop = main_genericstandalone_rx_cdc_fifo_out_eop;
assign main_genericstandalone_rx_cdc_source_payload_data = main_genericstandalone_rx_cdc_fifo_out_payload_data;
assign main_genericstandalone_rx_cdc_source_payload_last_be = main_genericstandalone_rx_cdc_fifo_out_payload_last_be;
assign main_genericstandalone_rx_cdc_source_payload_error = main_genericstandalone_rx_cdc_fifo_out_payload_error;
assign main_genericstandalone_rx_cdc_asyncfifo_re = main_genericstandalone_rx_cdc_source_ack;
assign main_genericstandalone_rx_cdc_graycounter0_ce = (main_genericstandalone_rx_cdc_asyncfifo_writable & main_genericstandalone_rx_cdc_asyncfifo_we);
assign main_genericstandalone_rx_cdc_graycounter1_ce = (main_genericstandalone_rx_cdc_asyncfifo_readable & main_genericstandalone_rx_cdc_asyncfifo_re);
assign main_genericstandalone_rx_cdc_asyncfifo_writable = (((main_genericstandalone_rx_cdc_graycounter0_q[6] == main_genericstandalone_rx_cdc_consume_wdomain[6]) | (main_genericstandalone_rx_cdc_graycounter0_q[5] == main_genericstandalone_rx_cdc_consume_wdomain[5])) | (main_genericstandalone_rx_cdc_graycounter0_q[4:0] != main_genericstandalone_rx_cdc_consume_wdomain[4:0]));
assign main_genericstandalone_rx_cdc_asyncfifo_readable = (main_genericstandalone_rx_cdc_graycounter1_q != main_genericstandalone_rx_cdc_produce_rdomain);
assign main_genericstandalone_rx_cdc_wrport_adr = main_genericstandalone_rx_cdc_graycounter0_q_binary[5:0];
assign main_genericstandalone_rx_cdc_wrport_dat_w = main_genericstandalone_rx_cdc_asyncfifo_din;
assign main_genericstandalone_rx_cdc_wrport_we = main_genericstandalone_rx_cdc_graycounter0_ce;
assign main_genericstandalone_rx_cdc_rdport_adr = main_genericstandalone_rx_cdc_graycounter1_q_next_binary[5:0];
assign main_genericstandalone_rx_cdc_asyncfifo_dout = main_genericstandalone_rx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_55;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_genericstandalone_rx_cdc_graycounter0_ce) begin
		main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= (main_genericstandalone_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_genericstandalone_rx_cdc_graycounter0_q_next_binary <= main_genericstandalone_rx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_55 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_cdc_graycounter0_q_next = (main_genericstandalone_rx_cdc_graycounter0_q_next_binary ^ main_genericstandalone_rx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_56;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_genericstandalone_rx_cdc_graycounter1_ce) begin
		main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= (main_genericstandalone_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_genericstandalone_rx_cdc_graycounter1_q_next_binary <= main_genericstandalone_rx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_56 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_rx_cdc_graycounter1_q_next = (main_genericstandalone_rx_cdc_graycounter1_q_next_binary ^ main_genericstandalone_rx_cdc_graycounter1_q_next_binary[6:1]);
assign main_genericstandalone_writer_sink_sink_stb = main_genericstandalone_sink_stb;
assign main_genericstandalone_sink_ack = main_genericstandalone_writer_sink_sink_ack;
assign main_genericstandalone_writer_sink_sink_eop = main_genericstandalone_sink_eop;
assign main_genericstandalone_writer_sink_sink_payload_data = main_genericstandalone_sink_payload_data;
assign main_genericstandalone_writer_sink_sink_payload_last_be = main_genericstandalone_sink_payload_last_be;
assign main_genericstandalone_writer_sink_sink_payload_error = main_genericstandalone_sink_payload_error;
assign main_genericstandalone_source_stb = main_genericstandalone_reader_source_source_stb;
assign main_genericstandalone_reader_source_source_ack = main_genericstandalone_source_ack;
assign main_genericstandalone_source_eop = main_genericstandalone_reader_source_source_eop;
assign main_genericstandalone_source_payload_data = main_genericstandalone_reader_source_source_payload_data;
assign main_genericstandalone_source_payload_last_be = main_genericstandalone_reader_source_source_payload_last_be;
assign main_genericstandalone_source_payload_error = main_genericstandalone_reader_source_source_payload_error;

// synthesis translate_off
reg dummy_d_57;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_writer_increment <= 3'd0;
	if (main_genericstandalone_writer_sink_sink_payload_last_be[3]) begin
		main_genericstandalone_writer_increment <= 1'd1;
	end else begin
		if (main_genericstandalone_writer_sink_sink_payload_last_be[2]) begin
			main_genericstandalone_writer_increment <= 2'd2;
		end else begin
			if (main_genericstandalone_writer_sink_sink_payload_last_be[1]) begin
				main_genericstandalone_writer_increment <= 2'd3;
			end else begin
				main_genericstandalone_writer_increment <= 3'd4;
			end
		end
	end
// synthesis translate_off
	dummy_d_57 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_writer_fifo_sink_payload_slot = main_genericstandalone_writer_slot;
assign main_genericstandalone_writer_fifo_sink_payload_length = main_genericstandalone_writer_counter;
assign main_genericstandalone_writer_fifo_source_ack = main_genericstandalone_writer_available_clear;
assign main_genericstandalone_writer_available_trigger = main_genericstandalone_writer_fifo_source_stb;
assign main_genericstandalone_writer_slot_status = main_genericstandalone_writer_fifo_source_payload_slot;
assign main_genericstandalone_writer_length_status = main_genericstandalone_writer_fifo_source_payload_length;

// synthesis translate_off
reg dummy_d_58;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_writer_memory0_adr <= 9'd0;
	main_genericstandalone_writer_memory0_we <= 1'd0;
	main_genericstandalone_writer_memory0_dat_w <= 32'd0;
	main_genericstandalone_writer_memory1_adr <= 9'd0;
	main_genericstandalone_writer_memory1_we <= 1'd0;
	main_genericstandalone_writer_memory1_dat_w <= 32'd0;
	main_genericstandalone_writer_memory2_adr <= 9'd0;
	main_genericstandalone_writer_memory2_we <= 1'd0;
	main_genericstandalone_writer_memory2_dat_w <= 32'd0;
	main_genericstandalone_writer_memory3_adr <= 9'd0;
	main_genericstandalone_writer_memory3_we <= 1'd0;
	main_genericstandalone_writer_memory3_dat_w <= 32'd0;
	case (main_genericstandalone_writer_slot)
		1'd0: begin
			main_genericstandalone_writer_memory0_adr <= main_genericstandalone_writer_counter[31:2];
			main_genericstandalone_writer_memory0_dat_w <= main_genericstandalone_writer_sink_sink_payload_data;
			if ((main_genericstandalone_writer_sink_sink_stb & main_genericstandalone_writer_ongoing)) begin
				main_genericstandalone_writer_memory0_we <= 4'd15;
			end
		end
		1'd1: begin
			main_genericstandalone_writer_memory1_adr <= main_genericstandalone_writer_counter[31:2];
			main_genericstandalone_writer_memory1_dat_w <= main_genericstandalone_writer_sink_sink_payload_data;
			if ((main_genericstandalone_writer_sink_sink_stb & main_genericstandalone_writer_ongoing)) begin
				main_genericstandalone_writer_memory1_we <= 4'd15;
			end
		end
		2'd2: begin
			main_genericstandalone_writer_memory2_adr <= main_genericstandalone_writer_counter[31:2];
			main_genericstandalone_writer_memory2_dat_w <= main_genericstandalone_writer_sink_sink_payload_data;
			if ((main_genericstandalone_writer_sink_sink_stb & main_genericstandalone_writer_ongoing)) begin
				main_genericstandalone_writer_memory2_we <= 4'd15;
			end
		end
		2'd3: begin
			main_genericstandalone_writer_memory3_adr <= main_genericstandalone_writer_counter[31:2];
			main_genericstandalone_writer_memory3_dat_w <= main_genericstandalone_writer_sink_sink_payload_data;
			if ((main_genericstandalone_writer_sink_sink_stb & main_genericstandalone_writer_ongoing)) begin
				main_genericstandalone_writer_memory3_we <= 4'd15;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_58 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_writer_status_w = main_genericstandalone_writer_available_status;

// synthesis translate_off
reg dummy_d_59;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_writer_available_clear <= 1'd0;
	if ((main_genericstandalone_writer_pending_re & main_genericstandalone_writer_pending_r)) begin
		main_genericstandalone_writer_available_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_59 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_writer_pending_w = main_genericstandalone_writer_available_pending;
assign main_genericstandalone_writer_irq = (main_genericstandalone_writer_pending_w & main_genericstandalone_writer_storage);
assign main_genericstandalone_writer_available_status = main_genericstandalone_writer_available_trigger;
assign main_genericstandalone_writer_available_pending = main_genericstandalone_writer_available_trigger;
assign main_genericstandalone_writer_fifo_syncfifo_din = {main_genericstandalone_writer_fifo_fifo_in_eop, main_genericstandalone_writer_fifo_fifo_in_payload_length, main_genericstandalone_writer_fifo_fifo_in_payload_slot};
assign {main_genericstandalone_writer_fifo_fifo_out_eop, main_genericstandalone_writer_fifo_fifo_out_payload_length, main_genericstandalone_writer_fifo_fifo_out_payload_slot} = main_genericstandalone_writer_fifo_syncfifo_dout;
assign main_genericstandalone_writer_fifo_sink_ack = main_genericstandalone_writer_fifo_syncfifo_writable;
assign main_genericstandalone_writer_fifo_syncfifo_we = main_genericstandalone_writer_fifo_sink_stb;
assign main_genericstandalone_writer_fifo_fifo_in_eop = main_genericstandalone_writer_fifo_sink_eop;
assign main_genericstandalone_writer_fifo_fifo_in_payload_slot = main_genericstandalone_writer_fifo_sink_payload_slot;
assign main_genericstandalone_writer_fifo_fifo_in_payload_length = main_genericstandalone_writer_fifo_sink_payload_length;
assign main_genericstandalone_writer_fifo_source_stb = main_genericstandalone_writer_fifo_syncfifo_readable;
assign main_genericstandalone_writer_fifo_source_eop = main_genericstandalone_writer_fifo_fifo_out_eop;
assign main_genericstandalone_writer_fifo_source_payload_slot = main_genericstandalone_writer_fifo_fifo_out_payload_slot;
assign main_genericstandalone_writer_fifo_source_payload_length = main_genericstandalone_writer_fifo_fifo_out_payload_length;
assign main_genericstandalone_writer_fifo_syncfifo_re = main_genericstandalone_writer_fifo_source_ack;

// synthesis translate_off
reg dummy_d_60;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_writer_fifo_wrport_adr <= 2'd0;
	if (main_genericstandalone_writer_fifo_replace) begin
		main_genericstandalone_writer_fifo_wrport_adr <= (main_genericstandalone_writer_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_writer_fifo_wrport_adr <= main_genericstandalone_writer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_60 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_writer_fifo_wrport_dat_w = main_genericstandalone_writer_fifo_syncfifo_din;
assign main_genericstandalone_writer_fifo_wrport_we = (main_genericstandalone_writer_fifo_syncfifo_we & (main_genericstandalone_writer_fifo_syncfifo_writable | main_genericstandalone_writer_fifo_replace));
assign main_genericstandalone_writer_fifo_do_read = (main_genericstandalone_writer_fifo_syncfifo_readable & main_genericstandalone_writer_fifo_syncfifo_re);
assign main_genericstandalone_writer_fifo_rdport_adr = main_genericstandalone_writer_fifo_consume;
assign main_genericstandalone_writer_fifo_syncfifo_dout = main_genericstandalone_writer_fifo_rdport_dat_r;
assign main_genericstandalone_writer_fifo_syncfifo_writable = (main_genericstandalone_writer_fifo_level != 3'd4);
assign main_genericstandalone_writer_fifo_syncfifo_readable = (main_genericstandalone_writer_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_61;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_writer_counter_reset <= 1'd0;
	main_genericstandalone_writer_counter_ce <= 1'd0;
	main_genericstandalone_writer_slot_ce <= 1'd0;
	main_genericstandalone_writer_ongoing <= 1'd0;
	main_genericstandalone_writer_fifo_sink_stb <= 1'd0;
	builder_liteethmacsramwriter_next_state <= 2'd0;
	main_genericstandalone_writer_errors_status_next_value <= 32'd0;
	main_genericstandalone_writer_errors_status_next_value_ce <= 1'd0;
	builder_liteethmacsramwriter_next_state <= builder_liteethmacsramwriter_state;
	case (builder_liteethmacsramwriter_state)
		1'd1: begin
			if (main_genericstandalone_writer_sink_sink_stb) begin
				if ((main_genericstandalone_writer_counter == 11'd1530)) begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end else begin
					main_genericstandalone_writer_counter_ce <= 1'd1;
					main_genericstandalone_writer_ongoing <= 1'd1;
				end
				if (main_genericstandalone_writer_sink_sink_eop) begin
					if (((main_genericstandalone_writer_sink_sink_payload_error & main_genericstandalone_writer_sink_sink_payload_last_be) != 1'd0)) begin
						main_genericstandalone_writer_counter_reset <= 1'd1;
						builder_liteethmacsramwriter_next_state <= 1'd0;
					end else begin
						builder_liteethmacsramwriter_next_state <= 2'd3;
					end
				end
			end
		end
		2'd2: begin
			main_genericstandalone_writer_counter_reset <= 1'd1;
			if ((main_genericstandalone_writer_sink_sink_stb & main_genericstandalone_writer_sink_sink_eop)) begin
				main_genericstandalone_writer_errors_status_next_value <= (main_genericstandalone_writer_errors_status + 1'd1);
				main_genericstandalone_writer_errors_status_next_value_ce <= 1'd1;
				builder_liteethmacsramwriter_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_genericstandalone_writer_counter_reset <= 1'd1;
			main_genericstandalone_writer_slot_ce <= 1'd1;
			main_genericstandalone_writer_fifo_sink_stb <= 1'd1;
			builder_liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (main_genericstandalone_writer_sink_sink_stb) begin
				if (main_genericstandalone_writer_fifo_sink_ack) begin
					main_genericstandalone_writer_ongoing <= 1'd1;
					main_genericstandalone_writer_counter_ce <= 1'd1;
					builder_liteethmacsramwriter_next_state <= 1'd1;
				end else begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_61 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_reader_fifo_sink_stb = main_genericstandalone_reader_start_re;
assign main_genericstandalone_reader_fifo_sink_payload_slot = main_genericstandalone_reader_slot_storage;
assign main_genericstandalone_reader_fifo_sink_payload_length = main_genericstandalone_reader_length_storage;
assign main_genericstandalone_reader_ready_status = main_genericstandalone_reader_fifo_sink_ack;

// synthesis translate_off
reg dummy_d_62;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_reader_source_source_payload_last_be <= 4'd0;
	if (main_genericstandalone_reader_last) begin
		if ((main_genericstandalone_reader_fifo_source_payload_length[1:0] == 2'd3)) begin
			main_genericstandalone_reader_source_source_payload_last_be <= 2'd2;
		end else begin
			if ((main_genericstandalone_reader_fifo_source_payload_length[1:0] == 2'd2)) begin
				main_genericstandalone_reader_source_source_payload_last_be <= 3'd4;
			end else begin
				if ((main_genericstandalone_reader_fifo_source_payload_length[1:0] == 1'd1)) begin
					main_genericstandalone_reader_source_source_payload_last_be <= 4'd8;
				end else begin
					main_genericstandalone_reader_source_source_payload_last_be <= 1'd1;
				end
			end
		end
	end
// synthesis translate_off
	dummy_d_62 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_reader_last = ((main_genericstandalone_reader_counter + 3'd4) >= main_genericstandalone_reader_fifo_source_payload_length);
assign main_genericstandalone_reader_memory0_adr = main_genericstandalone_reader_counter[10:2];
assign main_genericstandalone_reader_memory1_adr = main_genericstandalone_reader_counter[10:2];
assign main_genericstandalone_reader_memory2_adr = main_genericstandalone_reader_counter[10:2];
assign main_genericstandalone_reader_memory3_adr = main_genericstandalone_reader_counter[10:2];

// synthesis translate_off
reg dummy_d_63;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_reader_source_source_payload_data <= 32'd0;
	case (main_genericstandalone_reader_fifo_source_payload_slot)
		1'd0: begin
			main_genericstandalone_reader_source_source_payload_data <= main_genericstandalone_reader_memory0_dat_r;
		end
		1'd1: begin
			main_genericstandalone_reader_source_source_payload_data <= main_genericstandalone_reader_memory1_dat_r;
		end
		2'd2: begin
			main_genericstandalone_reader_source_source_payload_data <= main_genericstandalone_reader_memory2_dat_r;
		end
		2'd3: begin
			main_genericstandalone_reader_source_source_payload_data <= main_genericstandalone_reader_memory3_dat_r;
		end
	endcase
// synthesis translate_off
	dummy_d_63 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_reader_eventmanager_status_w = main_genericstandalone_reader_done_status;

// synthesis translate_off
reg dummy_d_64;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_reader_done_clear <= 1'd0;
	if ((main_genericstandalone_reader_eventmanager_pending_re & main_genericstandalone_reader_eventmanager_pending_r)) begin
		main_genericstandalone_reader_done_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_64 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_reader_eventmanager_pending_w = main_genericstandalone_reader_done_pending;
assign main_genericstandalone_reader_irq = (main_genericstandalone_reader_eventmanager_pending_w & main_genericstandalone_reader_eventmanager_storage);
assign main_genericstandalone_reader_done_status = 1'd0;
assign main_genericstandalone_reader_fifo_syncfifo_din = {main_genericstandalone_reader_fifo_fifo_in_eop, main_genericstandalone_reader_fifo_fifo_in_payload_length, main_genericstandalone_reader_fifo_fifo_in_payload_slot};
assign {main_genericstandalone_reader_fifo_fifo_out_eop, main_genericstandalone_reader_fifo_fifo_out_payload_length, main_genericstandalone_reader_fifo_fifo_out_payload_slot} = main_genericstandalone_reader_fifo_syncfifo_dout;
assign main_genericstandalone_reader_fifo_sink_ack = main_genericstandalone_reader_fifo_syncfifo_writable;
assign main_genericstandalone_reader_fifo_syncfifo_we = main_genericstandalone_reader_fifo_sink_stb;
assign main_genericstandalone_reader_fifo_fifo_in_eop = main_genericstandalone_reader_fifo_sink_eop;
assign main_genericstandalone_reader_fifo_fifo_in_payload_slot = main_genericstandalone_reader_fifo_sink_payload_slot;
assign main_genericstandalone_reader_fifo_fifo_in_payload_length = main_genericstandalone_reader_fifo_sink_payload_length;
assign main_genericstandalone_reader_fifo_source_stb = main_genericstandalone_reader_fifo_syncfifo_readable;
assign main_genericstandalone_reader_fifo_source_eop = main_genericstandalone_reader_fifo_fifo_out_eop;
assign main_genericstandalone_reader_fifo_source_payload_slot = main_genericstandalone_reader_fifo_fifo_out_payload_slot;
assign main_genericstandalone_reader_fifo_source_payload_length = main_genericstandalone_reader_fifo_fifo_out_payload_length;
assign main_genericstandalone_reader_fifo_syncfifo_re = main_genericstandalone_reader_fifo_source_ack;

// synthesis translate_off
reg dummy_d_65;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_reader_fifo_wrport_adr <= 2'd0;
	if (main_genericstandalone_reader_fifo_replace) begin
		main_genericstandalone_reader_fifo_wrport_adr <= (main_genericstandalone_reader_fifo_produce - 1'd1);
	end else begin
		main_genericstandalone_reader_fifo_wrport_adr <= main_genericstandalone_reader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_65 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_reader_fifo_wrport_dat_w = main_genericstandalone_reader_fifo_syncfifo_din;
assign main_genericstandalone_reader_fifo_wrport_we = (main_genericstandalone_reader_fifo_syncfifo_we & (main_genericstandalone_reader_fifo_syncfifo_writable | main_genericstandalone_reader_fifo_replace));
assign main_genericstandalone_reader_fifo_do_read = (main_genericstandalone_reader_fifo_syncfifo_readable & main_genericstandalone_reader_fifo_syncfifo_re);
assign main_genericstandalone_reader_fifo_rdport_adr = main_genericstandalone_reader_fifo_consume;
assign main_genericstandalone_reader_fifo_syncfifo_dout = main_genericstandalone_reader_fifo_rdport_dat_r;
assign main_genericstandalone_reader_fifo_syncfifo_writable = (main_genericstandalone_reader_fifo_level != 3'd4);
assign main_genericstandalone_reader_fifo_syncfifo_readable = (main_genericstandalone_reader_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_66;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_reader_source_source_stb <= 1'd0;
	main_genericstandalone_reader_source_source_eop <= 1'd0;
	main_genericstandalone_reader_done_trigger <= 1'd0;
	main_genericstandalone_reader_fifo_source_ack <= 1'd0;
	main_genericstandalone_reader_counter_reset <= 1'd0;
	main_genericstandalone_reader_counter_ce <= 1'd0;
	builder_liteethmacsramreader_next_state <= 2'd0;
	builder_liteethmacsramreader_next_state <= builder_liteethmacsramreader_state;
	case (builder_liteethmacsramreader_state)
		1'd1: begin
			if ((~main_genericstandalone_reader_last_d)) begin
				builder_liteethmacsramreader_next_state <= 2'd2;
			end else begin
				builder_liteethmacsramreader_next_state <= 2'd3;
			end
		end
		2'd2: begin
			main_genericstandalone_reader_source_source_stb <= 1'd1;
			main_genericstandalone_reader_source_source_eop <= main_genericstandalone_reader_last;
			if (main_genericstandalone_reader_source_source_ack) begin
				main_genericstandalone_reader_counter_ce <= (~main_genericstandalone_reader_last);
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
		2'd3: begin
			main_genericstandalone_reader_fifo_source_ack <= 1'd1;
			main_genericstandalone_reader_done_trigger <= 1'd1;
			builder_liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			main_genericstandalone_reader_counter_reset <= 1'd1;
			if (main_genericstandalone_reader_fifo_source_stb) begin
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_66 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_ev_irq = (main_genericstandalone_writer_irq | main_genericstandalone_reader_irq);
assign main_genericstandalone_sram0_adr0 = main_genericstandalone_sram0_bus_adr0[8:0];
assign main_genericstandalone_sram0_bus_dat_r0 = main_genericstandalone_sram0_dat_r0;
assign main_genericstandalone_sram1_adr0 = main_genericstandalone_sram1_bus_adr0[8:0];
assign main_genericstandalone_sram1_bus_dat_r0 = main_genericstandalone_sram1_dat_r0;
assign main_genericstandalone_sram2_adr0 = main_genericstandalone_sram2_bus_adr0[8:0];
assign main_genericstandalone_sram2_bus_dat_r0 = main_genericstandalone_sram2_dat_r0;
assign main_genericstandalone_sram3_adr0 = main_genericstandalone_sram3_bus_adr0[8:0];
assign main_genericstandalone_sram3_bus_dat_r0 = main_genericstandalone_sram3_dat_r0;

// synthesis translate_off
reg dummy_d_67;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram0_we <= 4'd0;
	main_genericstandalone_sram0_we[0] <= (((main_genericstandalone_sram0_bus_cyc1 & main_genericstandalone_sram0_bus_stb1) & main_genericstandalone_sram0_bus_we1) & main_genericstandalone_sram0_bus_sel1[0]);
	main_genericstandalone_sram0_we[1] <= (((main_genericstandalone_sram0_bus_cyc1 & main_genericstandalone_sram0_bus_stb1) & main_genericstandalone_sram0_bus_we1) & main_genericstandalone_sram0_bus_sel1[1]);
	main_genericstandalone_sram0_we[2] <= (((main_genericstandalone_sram0_bus_cyc1 & main_genericstandalone_sram0_bus_stb1) & main_genericstandalone_sram0_bus_we1) & main_genericstandalone_sram0_bus_sel1[2]);
	main_genericstandalone_sram0_we[3] <= (((main_genericstandalone_sram0_bus_cyc1 & main_genericstandalone_sram0_bus_stb1) & main_genericstandalone_sram0_bus_we1) & main_genericstandalone_sram0_bus_sel1[3]);
// synthesis translate_off
	dummy_d_67 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram0_adr1 = main_genericstandalone_sram0_bus_adr1[8:0];
assign main_genericstandalone_sram0_bus_dat_r1 = main_genericstandalone_sram0_dat_r1;
assign main_genericstandalone_sram0_dat_w = main_genericstandalone_sram0_bus_dat_w1;

// synthesis translate_off
reg dummy_d_68;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram1_we <= 4'd0;
	main_genericstandalone_sram1_we[0] <= (((main_genericstandalone_sram1_bus_cyc1 & main_genericstandalone_sram1_bus_stb1) & main_genericstandalone_sram1_bus_we1) & main_genericstandalone_sram1_bus_sel1[0]);
	main_genericstandalone_sram1_we[1] <= (((main_genericstandalone_sram1_bus_cyc1 & main_genericstandalone_sram1_bus_stb1) & main_genericstandalone_sram1_bus_we1) & main_genericstandalone_sram1_bus_sel1[1]);
	main_genericstandalone_sram1_we[2] <= (((main_genericstandalone_sram1_bus_cyc1 & main_genericstandalone_sram1_bus_stb1) & main_genericstandalone_sram1_bus_we1) & main_genericstandalone_sram1_bus_sel1[2]);
	main_genericstandalone_sram1_we[3] <= (((main_genericstandalone_sram1_bus_cyc1 & main_genericstandalone_sram1_bus_stb1) & main_genericstandalone_sram1_bus_we1) & main_genericstandalone_sram1_bus_sel1[3]);
// synthesis translate_off
	dummy_d_68 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram1_adr1 = main_genericstandalone_sram1_bus_adr1[8:0];
assign main_genericstandalone_sram1_bus_dat_r1 = main_genericstandalone_sram1_dat_r1;
assign main_genericstandalone_sram1_dat_w = main_genericstandalone_sram1_bus_dat_w1;

// synthesis translate_off
reg dummy_d_69;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram2_we <= 4'd0;
	main_genericstandalone_sram2_we[0] <= (((main_genericstandalone_sram2_bus_cyc1 & main_genericstandalone_sram2_bus_stb1) & main_genericstandalone_sram2_bus_we1) & main_genericstandalone_sram2_bus_sel1[0]);
	main_genericstandalone_sram2_we[1] <= (((main_genericstandalone_sram2_bus_cyc1 & main_genericstandalone_sram2_bus_stb1) & main_genericstandalone_sram2_bus_we1) & main_genericstandalone_sram2_bus_sel1[1]);
	main_genericstandalone_sram2_we[2] <= (((main_genericstandalone_sram2_bus_cyc1 & main_genericstandalone_sram2_bus_stb1) & main_genericstandalone_sram2_bus_we1) & main_genericstandalone_sram2_bus_sel1[2]);
	main_genericstandalone_sram2_we[3] <= (((main_genericstandalone_sram2_bus_cyc1 & main_genericstandalone_sram2_bus_stb1) & main_genericstandalone_sram2_bus_we1) & main_genericstandalone_sram2_bus_sel1[3]);
// synthesis translate_off
	dummy_d_69 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram2_adr1 = main_genericstandalone_sram2_bus_adr1[8:0];
assign main_genericstandalone_sram2_bus_dat_r1 = main_genericstandalone_sram2_dat_r1;
assign main_genericstandalone_sram2_dat_w = main_genericstandalone_sram2_bus_dat_w1;

// synthesis translate_off
reg dummy_d_70;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_sram3_we <= 4'd0;
	main_genericstandalone_sram3_we[0] <= (((main_genericstandalone_sram3_bus_cyc1 & main_genericstandalone_sram3_bus_stb1) & main_genericstandalone_sram3_bus_we1) & main_genericstandalone_sram3_bus_sel1[0]);
	main_genericstandalone_sram3_we[1] <= (((main_genericstandalone_sram3_bus_cyc1 & main_genericstandalone_sram3_bus_stb1) & main_genericstandalone_sram3_bus_we1) & main_genericstandalone_sram3_bus_sel1[1]);
	main_genericstandalone_sram3_we[2] <= (((main_genericstandalone_sram3_bus_cyc1 & main_genericstandalone_sram3_bus_stb1) & main_genericstandalone_sram3_bus_we1) & main_genericstandalone_sram3_bus_sel1[2]);
	main_genericstandalone_sram3_we[3] <= (((main_genericstandalone_sram3_bus_cyc1 & main_genericstandalone_sram3_bus_stb1) & main_genericstandalone_sram3_bus_we1) & main_genericstandalone_sram3_bus_sel1[3]);
// synthesis translate_off
	dummy_d_70 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram3_adr1 = main_genericstandalone_sram3_bus_adr1[8:0];
assign main_genericstandalone_sram3_bus_dat_r1 = main_genericstandalone_sram3_dat_r1;
assign main_genericstandalone_sram3_dat_w = main_genericstandalone_sram3_bus_dat_w1;

// synthesis translate_off
reg dummy_d_71;
// synthesis translate_on
always @(*) begin
	main_genericstandalone_slave_sel <= 8'd0;
	main_genericstandalone_slave_sel[0] <= (main_genericstandalone_bus_adr[11:9] == 1'd0);
	main_genericstandalone_slave_sel[1] <= (main_genericstandalone_bus_adr[11:9] == 1'd1);
	main_genericstandalone_slave_sel[2] <= (main_genericstandalone_bus_adr[11:9] == 2'd2);
	main_genericstandalone_slave_sel[3] <= (main_genericstandalone_bus_adr[11:9] == 2'd3);
	main_genericstandalone_slave_sel[4] <= (main_genericstandalone_bus_adr[11:9] == 3'd4);
	main_genericstandalone_slave_sel[5] <= (main_genericstandalone_bus_adr[11:9] == 3'd5);
	main_genericstandalone_slave_sel[6] <= (main_genericstandalone_bus_adr[11:9] == 3'd6);
	main_genericstandalone_slave_sel[7] <= (main_genericstandalone_bus_adr[11:9] == 3'd7);
// synthesis translate_off
	dummy_d_71 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_sram0_bus_adr0 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram0_bus_dat_w0 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram0_bus_sel0 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram0_bus_stb0 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram0_bus_we0 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram0_bus_cti0 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram0_bus_bte0 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram1_bus_adr0 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram1_bus_dat_w0 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram1_bus_sel0 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram1_bus_stb0 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram1_bus_we0 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram1_bus_cti0 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram1_bus_bte0 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram2_bus_adr0 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram2_bus_dat_w0 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram2_bus_sel0 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram2_bus_stb0 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram2_bus_we0 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram2_bus_cti0 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram2_bus_bte0 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram3_bus_adr0 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram3_bus_dat_w0 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram3_bus_sel0 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram3_bus_stb0 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram3_bus_we0 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram3_bus_cti0 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram3_bus_bte0 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram0_bus_adr1 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram0_bus_dat_w1 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram0_bus_sel1 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram0_bus_stb1 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram0_bus_we1 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram0_bus_cti1 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram0_bus_bte1 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram1_bus_adr1 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram1_bus_dat_w1 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram1_bus_sel1 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram1_bus_stb1 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram1_bus_we1 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram1_bus_cti1 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram1_bus_bte1 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram2_bus_adr1 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram2_bus_dat_w1 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram2_bus_sel1 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram2_bus_stb1 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram2_bus_we1 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram2_bus_cti1 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram2_bus_bte1 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram3_bus_adr1 = main_genericstandalone_bus_adr;
assign main_genericstandalone_sram3_bus_dat_w1 = main_genericstandalone_bus_dat_w;
assign main_genericstandalone_sram3_bus_sel1 = main_genericstandalone_bus_sel;
assign main_genericstandalone_sram3_bus_stb1 = main_genericstandalone_bus_stb;
assign main_genericstandalone_sram3_bus_we1 = main_genericstandalone_bus_we;
assign main_genericstandalone_sram3_bus_cti1 = main_genericstandalone_bus_cti;
assign main_genericstandalone_sram3_bus_bte1 = main_genericstandalone_bus_bte;
assign main_genericstandalone_sram0_bus_cyc0 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[0]);
assign main_genericstandalone_sram1_bus_cyc0 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[1]);
assign main_genericstandalone_sram2_bus_cyc0 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[2]);
assign main_genericstandalone_sram3_bus_cyc0 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[3]);
assign main_genericstandalone_sram0_bus_cyc1 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[4]);
assign main_genericstandalone_sram1_bus_cyc1 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[5]);
assign main_genericstandalone_sram2_bus_cyc1 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[6]);
assign main_genericstandalone_sram3_bus_cyc1 = (main_genericstandalone_bus_cyc & main_genericstandalone_slave_sel[7]);
assign main_genericstandalone_bus_ack = (((((((main_genericstandalone_sram0_bus_ack0 | main_genericstandalone_sram1_bus_ack0) | main_genericstandalone_sram2_bus_ack0) | main_genericstandalone_sram3_bus_ack0) | main_genericstandalone_sram0_bus_ack1) | main_genericstandalone_sram1_bus_ack1) | main_genericstandalone_sram2_bus_ack1) | main_genericstandalone_sram3_bus_ack1);
assign main_genericstandalone_bus_err = (((((((main_genericstandalone_sram0_bus_err0 | main_genericstandalone_sram1_bus_err0) | main_genericstandalone_sram2_bus_err0) | main_genericstandalone_sram3_bus_err0) | main_genericstandalone_sram0_bus_err1) | main_genericstandalone_sram1_bus_err1) | main_genericstandalone_sram2_bus_err1) | main_genericstandalone_sram3_bus_err1);
assign main_genericstandalone_bus_dat_r = (((((((({32{main_genericstandalone_slave_sel_r[0]}} & main_genericstandalone_sram0_bus_dat_r0) | ({32{main_genericstandalone_slave_sel_r[1]}} & main_genericstandalone_sram1_bus_dat_r0)) | ({32{main_genericstandalone_slave_sel_r[2]}} & main_genericstandalone_sram2_bus_dat_r0)) | ({32{main_genericstandalone_slave_sel_r[3]}} & main_genericstandalone_sram3_bus_dat_r0)) | ({32{main_genericstandalone_slave_sel_r[4]}} & main_genericstandalone_sram0_bus_dat_r1)) | ({32{main_genericstandalone_slave_sel_r[5]}} & main_genericstandalone_sram1_bus_dat_r1)) | ({32{main_genericstandalone_slave_sel_r[6]}} & main_genericstandalone_sram2_bus_dat_r1)) | ({32{main_genericstandalone_slave_sel_r[7]}} & main_genericstandalone_sram3_bus_dat_r1));
assign sys_kernel_clk = sys_clk;
assign sys_kernel_rst = main_genericstandalone_kernel_cpu_storage;
assign main_genericstandalone_kernel_cpu_ibus_adr = main_genericstandalone_kernel_cpu_i_adr_o[31:2];
assign main_genericstandalone_kernel_cpu_dbus_adr = main_genericstandalone_kernel_cpu_d_adr_o[31:2];
assign builder_shared_adr = builder_comb_rhs_array_muxed0;
assign builder_shared_dat_w = builder_comb_rhs_array_muxed1;
assign builder_shared_sel = builder_comb_rhs_array_muxed2;
assign builder_shared_cyc = builder_comb_rhs_array_muxed3;
assign builder_shared_stb = builder_comb_rhs_array_muxed4;
assign builder_shared_we = builder_comb_rhs_array_muxed5;
assign builder_shared_cti = builder_comb_rhs_array_muxed6;
assign builder_shared_bte = builder_comb_rhs_array_muxed7;
assign main_genericstandalone_kernel_cpu_ibus_dat_r = builder_shared_dat_r;
assign main_genericstandalone_kernel_cpu_dbus_dat_r = builder_shared_dat_r;
assign main_genericstandalone_kernel_cpu_ibus_ack = (builder_shared_ack & (builder_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_dbus_ack = (builder_shared_ack & (builder_grant == 1'd1));
assign main_genericstandalone_kernel_cpu_ibus_err = (builder_shared_err & (builder_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_dbus_err = (builder_shared_err & (builder_grant == 1'd1));
assign builder_request = {(main_genericstandalone_kernel_cpu_dbus_cyc & (~main_genericstandalone_kernel_cpu_dbus_ack)), (main_genericstandalone_kernel_cpu_ibus_cyc & (~main_genericstandalone_kernel_cpu_ibus_ack))};

// synthesis translate_off
reg dummy_d_72;
// synthesis translate_on
always @(*) begin
	builder_slave_sel <= 5'd0;
	builder_slave_sel[0] <= ((1'd1 & (~builder_shared_adr[27])) & builder_shared_adr[28]);
	builder_slave_sel[1] <= ((1'd1 & builder_shared_adr[27]) & builder_shared_adr[28]);
	builder_slave_sel[2] <= (((1'd1 & (~builder_shared_adr[26])) & (~builder_shared_adr[28])) & builder_shared_adr[27]);
	builder_slave_sel[3] <= (((1'd1 & (~builder_shared_adr[28])) & builder_shared_adr[26]) & builder_shared_adr[27]);
	builder_slave_sel[4] <= ((1'd1 & (~builder_shared_adr[27])) & (~builder_shared_adr[28]));
// synthesis translate_off
	dummy_d_72 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_kernel_cpu_wb_sdram_adr = builder_shared_adr;
assign main_genericstandalone_kernel_cpu_wb_sdram_dat_w = builder_shared_dat_w;
assign main_genericstandalone_kernel_cpu_wb_sdram_sel = builder_shared_sel;
assign main_genericstandalone_kernel_cpu_wb_sdram_stb = builder_shared_stb;
assign main_genericstandalone_kernel_cpu_wb_sdram_we = builder_shared_we;
assign main_genericstandalone_kernel_cpu_wb_sdram_cti = builder_shared_cti;
assign main_genericstandalone_kernel_cpu_wb_sdram_bte = builder_shared_bte;
assign main_genericstandalone_mailbox_i2_adr = builder_shared_adr;
assign main_genericstandalone_mailbox_i2_dat_w = builder_shared_dat_w;
assign main_genericstandalone_mailbox_i2_sel = builder_shared_sel;
assign main_genericstandalone_mailbox_i2_stb = builder_shared_stb;
assign main_genericstandalone_mailbox_i2_we = builder_shared_we;
assign main_genericstandalone_mailbox_i2_cti = builder_shared_cti;
assign main_genericstandalone_mailbox_i2_bte = builder_shared_bte;
assign main_genericstandalone_csrbank0_bus_adr = builder_shared_adr;
assign main_genericstandalone_csrbank0_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_csrbank0_bus_sel = builder_shared_sel;
assign main_genericstandalone_csrbank0_bus_stb = builder_shared_stb;
assign main_genericstandalone_csrbank0_bus_we = builder_shared_we;
assign main_genericstandalone_csrbank0_bus_cti = builder_shared_cti;
assign main_genericstandalone_csrbank0_bus_bte = builder_shared_bte;
assign main_genericstandalone_csrbank1_bus_adr = builder_shared_adr;
assign main_genericstandalone_csrbank1_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_csrbank1_bus_sel = builder_shared_sel;
assign main_genericstandalone_csrbank1_bus_stb = builder_shared_stb;
assign main_genericstandalone_csrbank1_bus_we = builder_shared_we;
assign main_genericstandalone_csrbank1_bus_cti = builder_shared_cti;
assign main_genericstandalone_csrbank1_bus_bte = builder_shared_bte;
assign main_genericstandalone_csrbank2_bus_adr = builder_shared_adr;
assign main_genericstandalone_csrbank2_bus_dat_w = builder_shared_dat_w;
assign main_genericstandalone_csrbank2_bus_sel = builder_shared_sel;
assign main_genericstandalone_csrbank2_bus_stb = builder_shared_stb;
assign main_genericstandalone_csrbank2_bus_we = builder_shared_we;
assign main_genericstandalone_csrbank2_bus_cti = builder_shared_cti;
assign main_genericstandalone_csrbank2_bus_bte = builder_shared_bte;
assign main_genericstandalone_kernel_cpu_wb_sdram_cyc = (builder_shared_cyc & builder_slave_sel[0]);
assign main_genericstandalone_mailbox_i2_cyc = (builder_shared_cyc & builder_slave_sel[1]);
assign main_genericstandalone_csrbank0_bus_cyc = (builder_shared_cyc & builder_slave_sel[2]);
assign main_genericstandalone_csrbank1_bus_cyc = (builder_shared_cyc & builder_slave_sel[3]);
assign main_genericstandalone_csrbank2_bus_cyc = (builder_shared_cyc & builder_slave_sel[4]);
assign builder_shared_ack = ((((main_genericstandalone_kernel_cpu_wb_sdram_ack | main_genericstandalone_mailbox_i2_ack) | main_genericstandalone_csrbank0_bus_ack) | main_genericstandalone_csrbank1_bus_ack) | main_genericstandalone_csrbank2_bus_ack);
assign builder_shared_err = ((((main_genericstandalone_kernel_cpu_wb_sdram_err | main_genericstandalone_mailbox_i2_err) | main_genericstandalone_csrbank0_bus_err) | main_genericstandalone_csrbank1_bus_err) | main_genericstandalone_csrbank2_bus_err);
assign builder_shared_dat_r = ((((({32{builder_slave_sel_r[0]}} & main_genericstandalone_kernel_cpu_wb_sdram_dat_r) | ({32{builder_slave_sel_r[1]}} & main_genericstandalone_mailbox_i2_dat_r)) | ({32{builder_slave_sel_r[2]}} & main_genericstandalone_csrbank0_bus_dat_r)) | ({32{builder_slave_sel_r[3]}} & main_genericstandalone_csrbank1_bus_dat_r)) | ({32{builder_slave_sel_r[4]}} & main_genericstandalone_csrbank2_bus_dat_r));
assign main_add_identifier_adr = main_add_identifier_storage;
assign main_add_identifier_status = main_add_identifier_dat_r;
assign {user_led} = main_leds_storage;
assign main_i2c_tstriple0_o = main_i2c_out_storage[0];
assign main_i2c_tstriple0_oe = main_i2c_oe_storage[0];

// synthesis translate_off
reg dummy_d_73;
// synthesis translate_on
always @(*) begin
	main_i2c_status0 <= 2'd0;
	main_i2c_status0[0] <= main_i2c_status1;
	main_i2c_status0[1] <= main_i2c_status2;
// synthesis translate_off
	dummy_d_73 <= dummy_s;
// synthesis translate_on
end
assign main_i2c_tstriple1_o = main_i2c_out_storage[1];
assign main_i2c_tstriple1_oe = main_i2c_oe_storage[1];
assign main_inout_8x0_inout_8x0_input_state = main_inout_8x0_serdes_i0[7];
assign main_inout_8x0_inout_8x0_i = (main_inout_8x0_serdes_i0 ^ {8{main_inout_8x0_inout_8x0_i_d}});
assign main_inout_8x0_serdes_i0 = main_inout_8x0_serdes_i1;
assign main_inout_8x0_serdes_t_in = (~main_inout_8x0_serdes_oe);
assign main_inout_8x0_serdes_o1 = main_inout_8x0_serdes_o0;
assign main_inout_8x0_serdes_pad_i1 = main_inout_8x0_serdes_pad_i0;
assign main_inout_8x0_serdes_pad_o0 = main_inout_8x0_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_74;
// synthesis translate_on
always @(*) begin
	main_inout_8x0_inout_8x0_o <= 3'd0;
	if (main_inout_8x0_inout_8x0_i[7]) begin
		main_inout_8x0_inout_8x0_o <= 3'd7;
	end
	if (main_inout_8x0_inout_8x0_i[6]) begin
		main_inout_8x0_inout_8x0_o <= 3'd6;
	end
	if (main_inout_8x0_inout_8x0_i[5]) begin
		main_inout_8x0_inout_8x0_o <= 3'd5;
	end
	if (main_inout_8x0_inout_8x0_i[4]) begin
		main_inout_8x0_inout_8x0_o <= 3'd4;
	end
	if (main_inout_8x0_inout_8x0_i[3]) begin
		main_inout_8x0_inout_8x0_o <= 2'd3;
	end
	if (main_inout_8x0_inout_8x0_i[2]) begin
		main_inout_8x0_inout_8x0_o <= 2'd2;
	end
	if (main_inout_8x0_inout_8x0_i[1]) begin
		main_inout_8x0_inout_8x0_o <= 1'd1;
	end
	if (main_inout_8x0_inout_8x0_i[0]) begin
		main_inout_8x0_inout_8x0_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_74 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x0_inout_8x0_n = (main_inout_8x0_inout_8x0_i == 1'd0);
assign main_inout_8x1_inout_8x1_input_state = main_inout_8x1_serdes_i0[7];
assign main_inout_8x1_inout_8x1_i = (main_inout_8x1_serdes_i0 ^ {8{main_inout_8x1_inout_8x1_i_d}});
assign main_inout_8x1_serdes_i0 = main_inout_8x1_serdes_i1;
assign main_inout_8x1_serdes_t_in = (~main_inout_8x1_serdes_oe);
assign main_inout_8x1_serdes_o1 = main_inout_8x1_serdes_o0;
assign main_inout_8x1_serdes_pad_i1 = main_inout_8x1_serdes_pad_i0;
assign main_inout_8x1_serdes_pad_o0 = main_inout_8x1_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_75;
// synthesis translate_on
always @(*) begin
	main_inout_8x1_inout_8x1_o <= 3'd0;
	if (main_inout_8x1_inout_8x1_i[7]) begin
		main_inout_8x1_inout_8x1_o <= 3'd7;
	end
	if (main_inout_8x1_inout_8x1_i[6]) begin
		main_inout_8x1_inout_8x1_o <= 3'd6;
	end
	if (main_inout_8x1_inout_8x1_i[5]) begin
		main_inout_8x1_inout_8x1_o <= 3'd5;
	end
	if (main_inout_8x1_inout_8x1_i[4]) begin
		main_inout_8x1_inout_8x1_o <= 3'd4;
	end
	if (main_inout_8x1_inout_8x1_i[3]) begin
		main_inout_8x1_inout_8x1_o <= 2'd3;
	end
	if (main_inout_8x1_inout_8x1_i[2]) begin
		main_inout_8x1_inout_8x1_o <= 2'd2;
	end
	if (main_inout_8x1_inout_8x1_i[1]) begin
		main_inout_8x1_inout_8x1_o <= 1'd1;
	end
	if (main_inout_8x1_inout_8x1_i[0]) begin
		main_inout_8x1_inout_8x1_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_75 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x1_inout_8x1_n = (main_inout_8x1_inout_8x1_i == 1'd0);
assign main_inout_8x2_inout_8x2_input_state = main_inout_8x2_serdes_i0[7];
assign main_inout_8x2_inout_8x2_i = (main_inout_8x2_serdes_i0 ^ {8{main_inout_8x2_inout_8x2_i_d}});
assign main_inout_8x2_serdes_i0 = main_inout_8x2_serdes_i1;
assign main_inout_8x2_serdes_t_in = (~main_inout_8x2_serdes_oe);
assign main_inout_8x2_serdes_o1 = main_inout_8x2_serdes_o0;
assign main_inout_8x2_serdes_pad_i1 = main_inout_8x2_serdes_pad_i0;
assign main_inout_8x2_serdes_pad_o0 = main_inout_8x2_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_76;
// synthesis translate_on
always @(*) begin
	main_inout_8x2_inout_8x2_o <= 3'd0;
	if (main_inout_8x2_inout_8x2_i[7]) begin
		main_inout_8x2_inout_8x2_o <= 3'd7;
	end
	if (main_inout_8x2_inout_8x2_i[6]) begin
		main_inout_8x2_inout_8x2_o <= 3'd6;
	end
	if (main_inout_8x2_inout_8x2_i[5]) begin
		main_inout_8x2_inout_8x2_o <= 3'd5;
	end
	if (main_inout_8x2_inout_8x2_i[4]) begin
		main_inout_8x2_inout_8x2_o <= 3'd4;
	end
	if (main_inout_8x2_inout_8x2_i[3]) begin
		main_inout_8x2_inout_8x2_o <= 2'd3;
	end
	if (main_inout_8x2_inout_8x2_i[2]) begin
		main_inout_8x2_inout_8x2_o <= 2'd2;
	end
	if (main_inout_8x2_inout_8x2_i[1]) begin
		main_inout_8x2_inout_8x2_o <= 1'd1;
	end
	if (main_inout_8x2_inout_8x2_i[0]) begin
		main_inout_8x2_inout_8x2_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_76 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x2_inout_8x2_n = (main_inout_8x2_inout_8x2_i == 1'd0);
assign main_inout_8x3_inout_8x3_input_state = main_inout_8x3_serdes_i0[7];
assign main_inout_8x3_inout_8x3_i = (main_inout_8x3_serdes_i0 ^ {8{main_inout_8x3_inout_8x3_i_d}});
assign main_inout_8x3_serdes_i0 = main_inout_8x3_serdes_i1;
assign main_inout_8x3_serdes_t_in = (~main_inout_8x3_serdes_oe);
assign main_inout_8x3_serdes_o1 = main_inout_8x3_serdes_o0;
assign main_inout_8x3_serdes_pad_i1 = main_inout_8x3_serdes_pad_i0;
assign main_inout_8x3_serdes_pad_o0 = main_inout_8x3_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_77;
// synthesis translate_on
always @(*) begin
	main_inout_8x3_inout_8x3_o <= 3'd0;
	if (main_inout_8x3_inout_8x3_i[7]) begin
		main_inout_8x3_inout_8x3_o <= 3'd7;
	end
	if (main_inout_8x3_inout_8x3_i[6]) begin
		main_inout_8x3_inout_8x3_o <= 3'd6;
	end
	if (main_inout_8x3_inout_8x3_i[5]) begin
		main_inout_8x3_inout_8x3_o <= 3'd5;
	end
	if (main_inout_8x3_inout_8x3_i[4]) begin
		main_inout_8x3_inout_8x3_o <= 3'd4;
	end
	if (main_inout_8x3_inout_8x3_i[3]) begin
		main_inout_8x3_inout_8x3_o <= 2'd3;
	end
	if (main_inout_8x3_inout_8x3_i[2]) begin
		main_inout_8x3_inout_8x3_o <= 2'd2;
	end
	if (main_inout_8x3_inout_8x3_i[1]) begin
		main_inout_8x3_inout_8x3_o <= 1'd1;
	end
	if (main_inout_8x3_inout_8x3_i[0]) begin
		main_inout_8x3_inout_8x3_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_77 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x3_inout_8x3_n = (main_inout_8x3_inout_8x3_i == 1'd0);
assign main_inout_8x4_inout_8x4_input_state = main_inout_8x4_serdes_i0[7];
assign main_inout_8x4_inout_8x4_i = (main_inout_8x4_serdes_i0 ^ {8{main_inout_8x4_inout_8x4_i_d}});
assign main_inout_8x4_serdes_i0 = main_inout_8x4_serdes_i1;
assign main_inout_8x4_serdes_t_in = (~main_inout_8x4_serdes_oe);
assign main_inout_8x4_serdes_o1 = main_inout_8x4_serdes_o0;
assign main_inout_8x4_serdes_pad_i1 = main_inout_8x4_serdes_pad_i0;
assign main_inout_8x4_serdes_pad_o0 = main_inout_8x4_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_78;
// synthesis translate_on
always @(*) begin
	main_inout_8x4_inout_8x4_o <= 3'd0;
	if (main_inout_8x4_inout_8x4_i[7]) begin
		main_inout_8x4_inout_8x4_o <= 3'd7;
	end
	if (main_inout_8x4_inout_8x4_i[6]) begin
		main_inout_8x4_inout_8x4_o <= 3'd6;
	end
	if (main_inout_8x4_inout_8x4_i[5]) begin
		main_inout_8x4_inout_8x4_o <= 3'd5;
	end
	if (main_inout_8x4_inout_8x4_i[4]) begin
		main_inout_8x4_inout_8x4_o <= 3'd4;
	end
	if (main_inout_8x4_inout_8x4_i[3]) begin
		main_inout_8x4_inout_8x4_o <= 2'd3;
	end
	if (main_inout_8x4_inout_8x4_i[2]) begin
		main_inout_8x4_inout_8x4_o <= 2'd2;
	end
	if (main_inout_8x4_inout_8x4_i[1]) begin
		main_inout_8x4_inout_8x4_o <= 1'd1;
	end
	if (main_inout_8x4_inout_8x4_i[0]) begin
		main_inout_8x4_inout_8x4_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_78 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x4_inout_8x4_n = (main_inout_8x4_inout_8x4_i == 1'd0);
assign main_inout_8x5_inout_8x5_input_state = main_inout_8x5_serdes_i0[7];
assign main_inout_8x5_inout_8x5_i = (main_inout_8x5_serdes_i0 ^ {8{main_inout_8x5_inout_8x5_i_d}});
assign main_inout_8x5_serdes_i0 = main_inout_8x5_serdes_i1;
assign main_inout_8x5_serdes_t_in = (~main_inout_8x5_serdes_oe);
assign main_inout_8x5_serdes_o1 = main_inout_8x5_serdes_o0;
assign main_inout_8x5_serdes_pad_i1 = main_inout_8x5_serdes_pad_i0;
assign main_inout_8x5_serdes_pad_o0 = main_inout_8x5_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_79;
// synthesis translate_on
always @(*) begin
	main_inout_8x5_inout_8x5_o <= 3'd0;
	if (main_inout_8x5_inout_8x5_i[7]) begin
		main_inout_8x5_inout_8x5_o <= 3'd7;
	end
	if (main_inout_8x5_inout_8x5_i[6]) begin
		main_inout_8x5_inout_8x5_o <= 3'd6;
	end
	if (main_inout_8x5_inout_8x5_i[5]) begin
		main_inout_8x5_inout_8x5_o <= 3'd5;
	end
	if (main_inout_8x5_inout_8x5_i[4]) begin
		main_inout_8x5_inout_8x5_o <= 3'd4;
	end
	if (main_inout_8x5_inout_8x5_i[3]) begin
		main_inout_8x5_inout_8x5_o <= 2'd3;
	end
	if (main_inout_8x5_inout_8x5_i[2]) begin
		main_inout_8x5_inout_8x5_o <= 2'd2;
	end
	if (main_inout_8x5_inout_8x5_i[1]) begin
		main_inout_8x5_inout_8x5_o <= 1'd1;
	end
	if (main_inout_8x5_inout_8x5_i[0]) begin
		main_inout_8x5_inout_8x5_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_79 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x5_inout_8x5_n = (main_inout_8x5_inout_8x5_i == 1'd0);
assign main_inout_8x6_inout_8x6_input_state = main_inout_8x6_serdes_i0[7];
assign main_inout_8x6_inout_8x6_i = (main_inout_8x6_serdes_i0 ^ {8{main_inout_8x6_inout_8x6_i_d}});
assign main_inout_8x6_serdes_i0 = main_inout_8x6_serdes_i1;
assign main_inout_8x6_serdes_t_in = (~main_inout_8x6_serdes_oe);
assign main_inout_8x6_serdes_o1 = main_inout_8x6_serdes_o0;
assign main_inout_8x6_serdes_pad_i1 = main_inout_8x6_serdes_pad_i0;
assign main_inout_8x6_serdes_pad_o0 = main_inout_8x6_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_80;
// synthesis translate_on
always @(*) begin
	main_inout_8x6_inout_8x6_o <= 3'd0;
	if (main_inout_8x6_inout_8x6_i[7]) begin
		main_inout_8x6_inout_8x6_o <= 3'd7;
	end
	if (main_inout_8x6_inout_8x6_i[6]) begin
		main_inout_8x6_inout_8x6_o <= 3'd6;
	end
	if (main_inout_8x6_inout_8x6_i[5]) begin
		main_inout_8x6_inout_8x6_o <= 3'd5;
	end
	if (main_inout_8x6_inout_8x6_i[4]) begin
		main_inout_8x6_inout_8x6_o <= 3'd4;
	end
	if (main_inout_8x6_inout_8x6_i[3]) begin
		main_inout_8x6_inout_8x6_o <= 2'd3;
	end
	if (main_inout_8x6_inout_8x6_i[2]) begin
		main_inout_8x6_inout_8x6_o <= 2'd2;
	end
	if (main_inout_8x6_inout_8x6_i[1]) begin
		main_inout_8x6_inout_8x6_o <= 1'd1;
	end
	if (main_inout_8x6_inout_8x6_i[0]) begin
		main_inout_8x6_inout_8x6_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_80 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x6_inout_8x6_n = (main_inout_8x6_inout_8x6_i == 1'd0);
assign main_inout_8x7_inout_8x7_input_state = main_inout_8x7_serdes_i0[7];
assign main_inout_8x7_inout_8x7_i = (main_inout_8x7_serdes_i0 ^ {8{main_inout_8x7_inout_8x7_i_d}});
assign main_inout_8x7_serdes_i0 = main_inout_8x7_serdes_i1;
assign main_inout_8x7_serdes_t_in = (~main_inout_8x7_serdes_oe);
assign main_inout_8x7_serdes_o1 = main_inout_8x7_serdes_o0;
assign main_inout_8x7_serdes_pad_i1 = main_inout_8x7_serdes_pad_i0;
assign main_inout_8x7_serdes_pad_o0 = main_inout_8x7_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_81;
// synthesis translate_on
always @(*) begin
	main_inout_8x7_inout_8x7_o <= 3'd0;
	if (main_inout_8x7_inout_8x7_i[7]) begin
		main_inout_8x7_inout_8x7_o <= 3'd7;
	end
	if (main_inout_8x7_inout_8x7_i[6]) begin
		main_inout_8x7_inout_8x7_o <= 3'd6;
	end
	if (main_inout_8x7_inout_8x7_i[5]) begin
		main_inout_8x7_inout_8x7_o <= 3'd5;
	end
	if (main_inout_8x7_inout_8x7_i[4]) begin
		main_inout_8x7_inout_8x7_o <= 3'd4;
	end
	if (main_inout_8x7_inout_8x7_i[3]) begin
		main_inout_8x7_inout_8x7_o <= 2'd3;
	end
	if (main_inout_8x7_inout_8x7_i[2]) begin
		main_inout_8x7_inout_8x7_o <= 2'd2;
	end
	if (main_inout_8x7_inout_8x7_i[1]) begin
		main_inout_8x7_inout_8x7_o <= 1'd1;
	end
	if (main_inout_8x7_inout_8x7_i[0]) begin
		main_inout_8x7_inout_8x7_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_81 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x7_inout_8x7_n = (main_inout_8x7_inout_8x7_i == 1'd0);
assign main_spimaster0_spimachine0_length = main_spimaster0_config_length;
assign main_spimaster0_spimachine0_end0 = main_spimaster0_config_end;
assign main_spimaster0_spimachine0_div = main_spimaster0_config_div;
assign main_spimaster0_spimachine0_clk_phase = main_spimaster0_config_clk_phase;
assign main_spimaster0_spimachine0_lsb_first = main_spimaster0_config_lsb_first;
assign main_spimaster0_interface_half_duplex = main_spimaster0_config_half_duplex;
assign main_spimaster0_interface_cs0 = main_spimaster0_config_cs;
assign main_spimaster0_interface_cs_polarity = {3{main_spimaster0_config_cs_polarity}};
assign main_spimaster0_interface_clk_polarity = main_spimaster0_config_clk_polarity;
assign main_spimaster0_interface_offline = main_spimaster0_config_offline;
assign main_spimaster0_interface_cs_next = main_spimaster0_spimachine0_cs_next;
assign main_spimaster0_interface_clk_next = main_spimaster0_spimachine0_clk_next;
assign main_spimaster0_interface_ce = main_spimaster0_spimachine0_ce;
assign main_spimaster0_interface_sample = main_spimaster0_spimachine0_sample;
assign main_spimaster0_spimachine0_sdi = main_spimaster0_interface_sdi;
assign main_spimaster0_interface_sdo = main_spimaster0_spimachine0_sdo;
assign main_spimaster0_spimachine0_load0 = ((main_spimaster0_ointerface0_stb & main_spimaster0_spimachine0_writable) & (~main_spimaster0_ointerface0_address));
assign main_spimaster0_spimachine0_pdo = main_spimaster0_ointerface0_data;
assign main_spimaster0_ointerface0_busy = (~main_spimaster0_spimachine0_writable);
assign main_spimaster0_iinterface0_stb = (main_spimaster0_spimachine0_readable & main_spimaster0_read);
assign main_spimaster0_iinterface0_data = main_spimaster0_spimachine0_pdi;
assign main_spimaster0_interface_sdi = (main_spimaster0_interface_half_duplex ? main_spimaster0_interface_mosi_reg : main_spimaster0_interface_miso_reg);
assign main_spimaster0_spimachine0_ce = (main_spimaster0_spimachine0_done & main_spimaster0_spimachine0_count);
assign main_spimaster0_spimachine0_pdi = (main_spimaster0_spimachine0_lsb_first ? {main_spimaster0_spimachine0_sdi, main_spimaster0_spimachine0_sr[31:1]} : {main_spimaster0_spimachine0_sr[30:0], main_spimaster0_spimachine0_sdi});
assign main_spimaster0_spimachine0_cnt_done = (main_spimaster0_spimachine0_cnt == 1'd0);
assign main_spimaster0_spimachine0_done = (main_spimaster0_spimachine0_cnt_done & (~main_spimaster0_spimachine0_do_extend));

// synthesis translate_off
reg dummy_d_82;
// synthesis translate_on
always @(*) begin
	main_spimaster0_spimachine0_clk_next <= 1'd0;
	main_spimaster0_spimachine0_cs_next <= 1'd0;
	main_spimaster0_spimachine0_idle <= 1'd0;
	main_spimaster0_spimachine0_readable <= 1'd0;
	main_spimaster0_spimachine0_writable <= 1'd0;
	main_spimaster0_spimachine0_load1 <= 1'd0;
	main_spimaster0_spimachine0_shift <= 1'd0;
	main_spimaster0_spimachine0_sample <= 1'd0;
	main_spimaster0_spimachine0_extend <= 1'd0;
	main_spimaster0_spimachine0_count <= 1'd0;
	builder_spimaster0_next_state <= 3'd0;
	builder_spimaster0_next_state <= builder_spimaster0_state;
	case (builder_spimaster0_state)
		1'd1: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_extend <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= 1'd1;
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= (~main_spimaster0_spimachine0_clk_phase);
			if (main_spimaster0_spimachine0_done) begin
				main_spimaster0_spimachine0_sample <= 1'd1;
				builder_spimaster0_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_extend <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= main_spimaster0_spimachine0_clk_phase;
			if (main_spimaster0_spimachine0_done) begin
				if ((main_spimaster0_spimachine0_n == 1'd0)) begin
					main_spimaster0_spimachine0_readable <= 1'd1;
					main_spimaster0_spimachine0_writable <= 1'd1;
					if (main_spimaster0_spimachine0_end1) begin
						main_spimaster0_spimachine0_clk_next <= 1'd0;
						main_spimaster0_spimachine0_writable <= 1'd0;
						if (main_spimaster0_spimachine0_clk_phase) begin
							main_spimaster0_spimachine0_cs_next <= 1'd0;
							builder_spimaster0_next_state <= 3'd5;
						end else begin
							builder_spimaster0_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster0_spimachine0_load0) begin
							main_spimaster0_spimachine0_load1 <= 1'd1;
							builder_spimaster0_next_state <= 2'd2;
						end else begin
							main_spimaster0_spimachine0_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster0_spimachine0_shift <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster0_spimachine0_count <= 1'd1;
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster0_spimachine0_idle <= 1'd1;
			main_spimaster0_spimachine0_writable <= 1'd1;
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			if (main_spimaster0_spimachine0_load0) begin
				main_spimaster0_spimachine0_count <= 1'd1;
				main_spimaster0_spimachine0_load1 <= 1'd1;
				if (main_spimaster0_spimachine0_clk_phase) begin
					builder_spimaster0_next_state <= 1'd1;
				end else begin
					main_spimaster0_spimachine0_extend <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_82 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster1_spimachine1_length = main_spimaster1_config_length;
assign main_spimaster1_spimachine1_end0 = main_spimaster1_config_end;
assign main_spimaster1_spimachine1_div = main_spimaster1_config_div;
assign main_spimaster1_spimachine1_clk_phase = main_spimaster1_config_clk_phase;
assign main_spimaster1_spimachine1_lsb_first = main_spimaster1_config_lsb_first;
assign main_spimaster1_interface_half_duplex = main_spimaster1_config_half_duplex;
assign main_spimaster1_interface_cs0 = main_spimaster1_config_cs;
assign main_spimaster1_interface_cs_polarity = {3{main_spimaster1_config_cs_polarity}};
assign main_spimaster1_interface_clk_polarity = main_spimaster1_config_clk_polarity;
assign main_spimaster1_interface_offline = main_spimaster1_config_offline;
assign main_spimaster1_interface_cs_next = main_spimaster1_spimachine1_cs_next;
assign main_spimaster1_interface_clk_next = main_spimaster1_spimachine1_clk_next;
assign main_spimaster1_interface_ce = main_spimaster1_spimachine1_ce;
assign main_spimaster1_interface_sample = main_spimaster1_spimachine1_sample;
assign main_spimaster1_spimachine1_sdi = main_spimaster1_interface_sdi;
assign main_spimaster1_interface_sdo = main_spimaster1_spimachine1_sdo;
assign main_spimaster1_spimachine1_load0 = ((main_spimaster1_ointerface1_stb & main_spimaster1_spimachine1_writable) & (~main_spimaster1_ointerface1_address));
assign main_spimaster1_spimachine1_pdo = main_spimaster1_ointerface1_data;
assign main_spimaster1_ointerface1_busy = (~main_spimaster1_spimachine1_writable);
assign main_spimaster1_iinterface1_stb = (main_spimaster1_spimachine1_readable & main_spimaster1_read);
assign main_spimaster1_iinterface1_data = main_spimaster1_spimachine1_pdi;
assign main_spimaster1_interface_sdi = (main_spimaster1_interface_half_duplex ? main_spimaster1_interface_mosi_reg : main_spimaster1_interface_miso_reg);
assign main_spimaster1_spimachine1_ce = (main_spimaster1_spimachine1_done & main_spimaster1_spimachine1_count);
assign main_spimaster1_spimachine1_pdi = (main_spimaster1_spimachine1_lsb_first ? {main_spimaster1_spimachine1_sdi, main_spimaster1_spimachine1_sr[31:1]} : {main_spimaster1_spimachine1_sr[30:0], main_spimaster1_spimachine1_sdi});
assign main_spimaster1_spimachine1_cnt_done = (main_spimaster1_spimachine1_cnt == 1'd0);
assign main_spimaster1_spimachine1_done = (main_spimaster1_spimachine1_cnt_done & (~main_spimaster1_spimachine1_do_extend));

// synthesis translate_off
reg dummy_d_83;
// synthesis translate_on
always @(*) begin
	main_spimaster1_spimachine1_clk_next <= 1'd0;
	main_spimaster1_spimachine1_cs_next <= 1'd0;
	main_spimaster1_spimachine1_idle <= 1'd0;
	main_spimaster1_spimachine1_readable <= 1'd0;
	main_spimaster1_spimachine1_writable <= 1'd0;
	main_spimaster1_spimachine1_load1 <= 1'd0;
	main_spimaster1_spimachine1_shift <= 1'd0;
	main_spimaster1_spimachine1_sample <= 1'd0;
	main_spimaster1_spimachine1_extend <= 1'd0;
	main_spimaster1_spimachine1_count <= 1'd0;
	builder_spimaster1_next_state <= 3'd0;
	builder_spimaster1_next_state <= builder_spimaster1_state;
	case (builder_spimaster1_state)
		1'd1: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_extend <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= 1'd1;
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= (~main_spimaster1_spimachine1_clk_phase);
			if (main_spimaster1_spimachine1_done) begin
				main_spimaster1_spimachine1_sample <= 1'd1;
				builder_spimaster1_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_extend <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= main_spimaster1_spimachine1_clk_phase;
			if (main_spimaster1_spimachine1_done) begin
				if ((main_spimaster1_spimachine1_n == 1'd0)) begin
					main_spimaster1_spimachine1_readable <= 1'd1;
					main_spimaster1_spimachine1_writable <= 1'd1;
					if (main_spimaster1_spimachine1_end1) begin
						main_spimaster1_spimachine1_clk_next <= 1'd0;
						main_spimaster1_spimachine1_writable <= 1'd0;
						if (main_spimaster1_spimachine1_clk_phase) begin
							main_spimaster1_spimachine1_cs_next <= 1'd0;
							builder_spimaster1_next_state <= 3'd5;
						end else begin
							builder_spimaster1_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster1_spimachine1_load0) begin
							main_spimaster1_spimachine1_load1 <= 1'd1;
							builder_spimaster1_next_state <= 2'd2;
						end else begin
							main_spimaster1_spimachine1_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster1_spimachine1_shift <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster1_spimachine1_count <= 1'd1;
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster1_spimachine1_idle <= 1'd1;
			main_spimaster1_spimachine1_writable <= 1'd1;
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			if (main_spimaster1_spimachine1_load0) begin
				main_spimaster1_spimachine1_count <= 1'd1;
				main_spimaster1_spimachine1_load1 <= 1'd1;
				if (main_spimaster1_spimachine1_clk_phase) begin
					builder_spimaster1_next_state <= 1'd1;
				end else begin
					main_spimaster1_spimachine1_extend <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_83 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster2_spimachine2_length = main_spimaster2_config_length;
assign main_spimaster2_spimachine2_end0 = main_spimaster2_config_end;
assign main_spimaster2_spimachine2_div = main_spimaster2_config_div;
assign main_spimaster2_spimachine2_clk_phase = main_spimaster2_config_clk_phase;
assign main_spimaster2_spimachine2_lsb_first = main_spimaster2_config_lsb_first;
assign main_spimaster2_interface_half_duplex = main_spimaster2_config_half_duplex;
assign main_spimaster2_interface_cs0 = main_spimaster2_config_cs;
assign main_spimaster2_interface_cs_polarity = {3{main_spimaster2_config_cs_polarity}};
assign main_spimaster2_interface_clk_polarity = main_spimaster2_config_clk_polarity;
assign main_spimaster2_interface_offline = main_spimaster2_config_offline;
assign main_spimaster2_interface_cs_next = main_spimaster2_spimachine2_cs_next;
assign main_spimaster2_interface_clk_next = main_spimaster2_spimachine2_clk_next;
assign main_spimaster2_interface_ce = main_spimaster2_spimachine2_ce;
assign main_spimaster2_interface_sample = main_spimaster2_spimachine2_sample;
assign main_spimaster2_spimachine2_sdi = main_spimaster2_interface_sdi;
assign main_spimaster2_interface_sdo = main_spimaster2_spimachine2_sdo;
assign main_spimaster2_spimachine2_load0 = ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable) & (~main_spimaster2_ointerface2_address));
assign main_spimaster2_spimachine2_pdo = main_spimaster2_ointerface2_data;
assign main_spimaster2_ointerface2_busy = (~main_spimaster2_spimachine2_writable);
assign main_spimaster2_iinterface2_stb = (main_spimaster2_spimachine2_readable & main_spimaster2_read);
assign main_spimaster2_iinterface2_data = main_spimaster2_spimachine2_pdi;
assign main_spimaster2_interface_sdi = (main_spimaster2_interface_half_duplex ? main_spimaster2_interface_mosi_reg : main_spimaster2_interface_miso_reg);
assign main_spimaster2_spimachine2_ce = (main_spimaster2_spimachine2_done & main_spimaster2_spimachine2_count);
assign main_spimaster2_spimachine2_pdi = (main_spimaster2_spimachine2_lsb_first ? {main_spimaster2_spimachine2_sdi, main_spimaster2_spimachine2_sr[31:1]} : {main_spimaster2_spimachine2_sr[30:0], main_spimaster2_spimachine2_sdi});
assign main_spimaster2_spimachine2_cnt_done = (main_spimaster2_spimachine2_cnt == 1'd0);
assign main_spimaster2_spimachine2_done = (main_spimaster2_spimachine2_cnt_done & (~main_spimaster2_spimachine2_do_extend));

// synthesis translate_off
reg dummy_d_84;
// synthesis translate_on
always @(*) begin
	main_spimaster2_spimachine2_clk_next <= 1'd0;
	main_spimaster2_spimachine2_cs_next <= 1'd0;
	main_spimaster2_spimachine2_idle <= 1'd0;
	main_spimaster2_spimachine2_readable <= 1'd0;
	main_spimaster2_spimachine2_writable <= 1'd0;
	main_spimaster2_spimachine2_load1 <= 1'd0;
	main_spimaster2_spimachine2_shift <= 1'd0;
	main_spimaster2_spimachine2_sample <= 1'd0;
	main_spimaster2_spimachine2_extend <= 1'd0;
	main_spimaster2_spimachine2_count <= 1'd0;
	builder_spimaster2_next_state <= 3'd0;
	builder_spimaster2_next_state <= builder_spimaster2_state;
	case (builder_spimaster2_state)
		1'd1: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= (~main_spimaster2_spimachine2_clk_phase);
			if (main_spimaster2_spimachine2_done) begin
				main_spimaster2_spimachine2_sample <= 1'd1;
				builder_spimaster2_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= main_spimaster2_spimachine2_clk_phase;
			if (main_spimaster2_spimachine2_done) begin
				if ((main_spimaster2_spimachine2_n == 1'd0)) begin
					main_spimaster2_spimachine2_readable <= 1'd1;
					main_spimaster2_spimachine2_writable <= 1'd1;
					if (main_spimaster2_spimachine2_end1) begin
						main_spimaster2_spimachine2_clk_next <= 1'd0;
						main_spimaster2_spimachine2_writable <= 1'd0;
						if (main_spimaster2_spimachine2_clk_phase) begin
							main_spimaster2_spimachine2_cs_next <= 1'd0;
							builder_spimaster2_next_state <= 3'd5;
						end else begin
							builder_spimaster2_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster2_spimachine2_load0) begin
							main_spimaster2_spimachine2_load1 <= 1'd1;
							builder_spimaster2_next_state <= 2'd2;
						end else begin
							main_spimaster2_spimachine2_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster2_spimachine2_shift <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster2_spimachine2_count <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster2_spimachine2_idle <= 1'd1;
			main_spimaster2_spimachine2_writable <= 1'd1;
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			if (main_spimaster2_spimachine2_load0) begin
				main_spimaster2_spimachine2_count <= 1'd1;
				main_spimaster2_spimachine2_load1 <= 1'd1;
				if (main_spimaster2_spimachine2_clk_phase) begin
					builder_spimaster2_next_state <= 1'd1;
				end else begin
					main_spimaster2_spimachine2_extend <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_84 <= dummy_s;
// synthesis translate_on
end
assign sfp_ctl_led_1 = main_output0_pad_o;
assign sfp_ctl_led_2 = main_output1_pad_o;
assign main_rtio_tsc_i = main_rtio_tsc_coarse_ts;
assign main_rtio_tsc_coarse_ts_sys = main_rtio_tsc_o;
assign main_rtio_tsc_full_ts = (main_rtio_tsc_coarse_ts <<< 2'd3);
assign main_rtio_tsc_full_ts_sys = (main_rtio_tsc_coarse_ts_sys <<< 2'd3);

// synthesis translate_off
reg dummy_d_85;
// synthesis translate_on
always @(*) begin
	main_rtio_tsc_value_sys <= 61'd0;
	main_rtio_tsc_value_sys[60] <= main_rtio_tsc_value_gray_sys[60];
	main_rtio_tsc_value_sys[59] <= (main_rtio_tsc_value_sys[60] ^ main_rtio_tsc_value_gray_sys[59]);
	main_rtio_tsc_value_sys[58] <= (main_rtio_tsc_value_sys[59] ^ main_rtio_tsc_value_gray_sys[58]);
	main_rtio_tsc_value_sys[57] <= (main_rtio_tsc_value_sys[58] ^ main_rtio_tsc_value_gray_sys[57]);
	main_rtio_tsc_value_sys[56] <= (main_rtio_tsc_value_sys[57] ^ main_rtio_tsc_value_gray_sys[56]);
	main_rtio_tsc_value_sys[55] <= (main_rtio_tsc_value_sys[56] ^ main_rtio_tsc_value_gray_sys[55]);
	main_rtio_tsc_value_sys[54] <= (main_rtio_tsc_value_sys[55] ^ main_rtio_tsc_value_gray_sys[54]);
	main_rtio_tsc_value_sys[53] <= (main_rtio_tsc_value_sys[54] ^ main_rtio_tsc_value_gray_sys[53]);
	main_rtio_tsc_value_sys[52] <= (main_rtio_tsc_value_sys[53] ^ main_rtio_tsc_value_gray_sys[52]);
	main_rtio_tsc_value_sys[51] <= (main_rtio_tsc_value_sys[52] ^ main_rtio_tsc_value_gray_sys[51]);
	main_rtio_tsc_value_sys[50] <= (main_rtio_tsc_value_sys[51] ^ main_rtio_tsc_value_gray_sys[50]);
	main_rtio_tsc_value_sys[49] <= (main_rtio_tsc_value_sys[50] ^ main_rtio_tsc_value_gray_sys[49]);
	main_rtio_tsc_value_sys[48] <= (main_rtio_tsc_value_sys[49] ^ main_rtio_tsc_value_gray_sys[48]);
	main_rtio_tsc_value_sys[47] <= (main_rtio_tsc_value_sys[48] ^ main_rtio_tsc_value_gray_sys[47]);
	main_rtio_tsc_value_sys[46] <= (main_rtio_tsc_value_sys[47] ^ main_rtio_tsc_value_gray_sys[46]);
	main_rtio_tsc_value_sys[45] <= (main_rtio_tsc_value_sys[46] ^ main_rtio_tsc_value_gray_sys[45]);
	main_rtio_tsc_value_sys[44] <= (main_rtio_tsc_value_sys[45] ^ main_rtio_tsc_value_gray_sys[44]);
	main_rtio_tsc_value_sys[43] <= (main_rtio_tsc_value_sys[44] ^ main_rtio_tsc_value_gray_sys[43]);
	main_rtio_tsc_value_sys[42] <= (main_rtio_tsc_value_sys[43] ^ main_rtio_tsc_value_gray_sys[42]);
	main_rtio_tsc_value_sys[41] <= (main_rtio_tsc_value_sys[42] ^ main_rtio_tsc_value_gray_sys[41]);
	main_rtio_tsc_value_sys[40] <= (main_rtio_tsc_value_sys[41] ^ main_rtio_tsc_value_gray_sys[40]);
	main_rtio_tsc_value_sys[39] <= (main_rtio_tsc_value_sys[40] ^ main_rtio_tsc_value_gray_sys[39]);
	main_rtio_tsc_value_sys[38] <= (main_rtio_tsc_value_sys[39] ^ main_rtio_tsc_value_gray_sys[38]);
	main_rtio_tsc_value_sys[37] <= (main_rtio_tsc_value_sys[38] ^ main_rtio_tsc_value_gray_sys[37]);
	main_rtio_tsc_value_sys[36] <= (main_rtio_tsc_value_sys[37] ^ main_rtio_tsc_value_gray_sys[36]);
	main_rtio_tsc_value_sys[35] <= (main_rtio_tsc_value_sys[36] ^ main_rtio_tsc_value_gray_sys[35]);
	main_rtio_tsc_value_sys[34] <= (main_rtio_tsc_value_sys[35] ^ main_rtio_tsc_value_gray_sys[34]);
	main_rtio_tsc_value_sys[33] <= (main_rtio_tsc_value_sys[34] ^ main_rtio_tsc_value_gray_sys[33]);
	main_rtio_tsc_value_sys[32] <= (main_rtio_tsc_value_sys[33] ^ main_rtio_tsc_value_gray_sys[32]);
	main_rtio_tsc_value_sys[31] <= (main_rtio_tsc_value_sys[32] ^ main_rtio_tsc_value_gray_sys[31]);
	main_rtio_tsc_value_sys[30] <= (main_rtio_tsc_value_sys[31] ^ main_rtio_tsc_value_gray_sys[30]);
	main_rtio_tsc_value_sys[29] <= (main_rtio_tsc_value_sys[30] ^ main_rtio_tsc_value_gray_sys[29]);
	main_rtio_tsc_value_sys[28] <= (main_rtio_tsc_value_sys[29] ^ main_rtio_tsc_value_gray_sys[28]);
	main_rtio_tsc_value_sys[27] <= (main_rtio_tsc_value_sys[28] ^ main_rtio_tsc_value_gray_sys[27]);
	main_rtio_tsc_value_sys[26] <= (main_rtio_tsc_value_sys[27] ^ main_rtio_tsc_value_gray_sys[26]);
	main_rtio_tsc_value_sys[25] <= (main_rtio_tsc_value_sys[26] ^ main_rtio_tsc_value_gray_sys[25]);
	main_rtio_tsc_value_sys[24] <= (main_rtio_tsc_value_sys[25] ^ main_rtio_tsc_value_gray_sys[24]);
	main_rtio_tsc_value_sys[23] <= (main_rtio_tsc_value_sys[24] ^ main_rtio_tsc_value_gray_sys[23]);
	main_rtio_tsc_value_sys[22] <= (main_rtio_tsc_value_sys[23] ^ main_rtio_tsc_value_gray_sys[22]);
	main_rtio_tsc_value_sys[21] <= (main_rtio_tsc_value_sys[22] ^ main_rtio_tsc_value_gray_sys[21]);
	main_rtio_tsc_value_sys[20] <= (main_rtio_tsc_value_sys[21] ^ main_rtio_tsc_value_gray_sys[20]);
	main_rtio_tsc_value_sys[19] <= (main_rtio_tsc_value_sys[20] ^ main_rtio_tsc_value_gray_sys[19]);
	main_rtio_tsc_value_sys[18] <= (main_rtio_tsc_value_sys[19] ^ main_rtio_tsc_value_gray_sys[18]);
	main_rtio_tsc_value_sys[17] <= (main_rtio_tsc_value_sys[18] ^ main_rtio_tsc_value_gray_sys[17]);
	main_rtio_tsc_value_sys[16] <= (main_rtio_tsc_value_sys[17] ^ main_rtio_tsc_value_gray_sys[16]);
	main_rtio_tsc_value_sys[15] <= (main_rtio_tsc_value_sys[16] ^ main_rtio_tsc_value_gray_sys[15]);
	main_rtio_tsc_value_sys[14] <= (main_rtio_tsc_value_sys[15] ^ main_rtio_tsc_value_gray_sys[14]);
	main_rtio_tsc_value_sys[13] <= (main_rtio_tsc_value_sys[14] ^ main_rtio_tsc_value_gray_sys[13]);
	main_rtio_tsc_value_sys[12] <= (main_rtio_tsc_value_sys[13] ^ main_rtio_tsc_value_gray_sys[12]);
	main_rtio_tsc_value_sys[11] <= (main_rtio_tsc_value_sys[12] ^ main_rtio_tsc_value_gray_sys[11]);
	main_rtio_tsc_value_sys[10] <= (main_rtio_tsc_value_sys[11] ^ main_rtio_tsc_value_gray_sys[10]);
	main_rtio_tsc_value_sys[9] <= (main_rtio_tsc_value_sys[10] ^ main_rtio_tsc_value_gray_sys[9]);
	main_rtio_tsc_value_sys[8] <= (main_rtio_tsc_value_sys[9] ^ main_rtio_tsc_value_gray_sys[8]);
	main_rtio_tsc_value_sys[7] <= (main_rtio_tsc_value_sys[8] ^ main_rtio_tsc_value_gray_sys[7]);
	main_rtio_tsc_value_sys[6] <= (main_rtio_tsc_value_sys[7] ^ main_rtio_tsc_value_gray_sys[6]);
	main_rtio_tsc_value_sys[5] <= (main_rtio_tsc_value_sys[6] ^ main_rtio_tsc_value_gray_sys[5]);
	main_rtio_tsc_value_sys[4] <= (main_rtio_tsc_value_sys[5] ^ main_rtio_tsc_value_gray_sys[4]);
	main_rtio_tsc_value_sys[3] <= (main_rtio_tsc_value_sys[4] ^ main_rtio_tsc_value_gray_sys[3]);
	main_rtio_tsc_value_sys[2] <= (main_rtio_tsc_value_sys[3] ^ main_rtio_tsc_value_gray_sys[2]);
	main_rtio_tsc_value_sys[1] <= (main_rtio_tsc_value_sys[2] ^ main_rtio_tsc_value_gray_sys[1]);
	main_rtio_tsc_value_sys[0] <= (main_rtio_tsc_value_sys[1] ^ main_rtio_tsc_value_gray_sys[0]);
// synthesis translate_off
	dummy_d_85 <= dummy_s;
// synthesis translate_on
end
assign rsys_clk = sys_clk;
assign rsys_rst = main_rtio_core_cmd_reset;
assign rio_clk = rtio_clk;
assign rio_phy_clk = rtio_clk;
assign main_rtio_core_outputs_gates_coarse_timestamp = main_rtio_tsc_coarse_ts;
assign main_rtio_core_async_error_w = {main_rtio_core_o_sequence_error, main_rtio_core_o_busy, main_rtio_core_o_collision};
assign main_rtio_core_o_collision_sync_i = main_rtio_core_outputs_collision;
assign main_rtio_core_o_collision_sync_data_i = main_rtio_core_outputs_collision_channel;
assign main_rtio_core_o_busy_sync_i = main_rtio_core_outputs_busy;
assign main_rtio_core_o_busy_sync_data_i = main_rtio_core_outputs_busy_channel;
assign main_rtio_core_outputs_record0_we = main_rtio_core_outputs_lanedistributor_record0_we;
assign main_rtio_core_outputs_lanedistributor_record0_writable = main_rtio_core_outputs_record0_writable;
assign main_rtio_core_outputs_record0_seqn0 = main_rtio_core_outputs_lanedistributor_record0_seqn;
assign main_rtio_core_outputs_record0_payload_channel0 = main_rtio_core_outputs_lanedistributor_record0_payload_channel;
assign main_rtio_core_outputs_record0_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
assign main_rtio_core_outputs_record0_payload_address0 = main_rtio_core_outputs_lanedistributor_record0_payload_address;
assign main_rtio_core_outputs_record0_payload_data0 = main_rtio_core_outputs_lanedistributor_record0_payload_data;
assign main_rtio_core_outputs_record1_we = main_rtio_core_outputs_lanedistributor_record1_we;
assign main_rtio_core_outputs_lanedistributor_record1_writable = main_rtio_core_outputs_record1_writable;
assign main_rtio_core_outputs_record1_seqn0 = main_rtio_core_outputs_lanedistributor_record1_seqn;
assign main_rtio_core_outputs_record1_payload_channel0 = main_rtio_core_outputs_lanedistributor_record1_payload_channel;
assign main_rtio_core_outputs_record1_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
assign main_rtio_core_outputs_record1_payload_address0 = main_rtio_core_outputs_lanedistributor_record1_payload_address;
assign main_rtio_core_outputs_record1_payload_data0 = main_rtio_core_outputs_lanedistributor_record1_payload_data;
assign main_rtio_core_outputs_record2_we = main_rtio_core_outputs_lanedistributor_record2_we;
assign main_rtio_core_outputs_lanedistributor_record2_writable = main_rtio_core_outputs_record2_writable;
assign main_rtio_core_outputs_record2_seqn0 = main_rtio_core_outputs_lanedistributor_record2_seqn;
assign main_rtio_core_outputs_record2_payload_channel0 = main_rtio_core_outputs_lanedistributor_record2_payload_channel;
assign main_rtio_core_outputs_record2_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
assign main_rtio_core_outputs_record2_payload_address0 = main_rtio_core_outputs_lanedistributor_record2_payload_address;
assign main_rtio_core_outputs_record2_payload_data0 = main_rtio_core_outputs_lanedistributor_record2_payload_data;
assign main_rtio_core_outputs_record3_we = main_rtio_core_outputs_lanedistributor_record3_we;
assign main_rtio_core_outputs_lanedistributor_record3_writable = main_rtio_core_outputs_record3_writable;
assign main_rtio_core_outputs_record3_seqn0 = main_rtio_core_outputs_lanedistributor_record3_seqn;
assign main_rtio_core_outputs_record3_payload_channel0 = main_rtio_core_outputs_lanedistributor_record3_payload_channel;
assign main_rtio_core_outputs_record3_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
assign main_rtio_core_outputs_record3_payload_address0 = main_rtio_core_outputs_lanedistributor_record3_payload_address;
assign main_rtio_core_outputs_record3_payload_data0 = main_rtio_core_outputs_lanedistributor_record3_payload_data;
assign main_rtio_core_outputs_record4_we = main_rtio_core_outputs_lanedistributor_record4_we;
assign main_rtio_core_outputs_lanedistributor_record4_writable = main_rtio_core_outputs_record4_writable;
assign main_rtio_core_outputs_record4_seqn0 = main_rtio_core_outputs_lanedistributor_record4_seqn;
assign main_rtio_core_outputs_record4_payload_channel0 = main_rtio_core_outputs_lanedistributor_record4_payload_channel;
assign main_rtio_core_outputs_record4_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
assign main_rtio_core_outputs_record4_payload_address0 = main_rtio_core_outputs_lanedistributor_record4_payload_address;
assign main_rtio_core_outputs_record4_payload_data0 = main_rtio_core_outputs_lanedistributor_record4_payload_data;
assign main_rtio_core_outputs_record5_we = main_rtio_core_outputs_lanedistributor_record5_we;
assign main_rtio_core_outputs_lanedistributor_record5_writable = main_rtio_core_outputs_record5_writable;
assign main_rtio_core_outputs_record5_seqn0 = main_rtio_core_outputs_lanedistributor_record5_seqn;
assign main_rtio_core_outputs_record5_payload_channel0 = main_rtio_core_outputs_lanedistributor_record5_payload_channel;
assign main_rtio_core_outputs_record5_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
assign main_rtio_core_outputs_record5_payload_address0 = main_rtio_core_outputs_lanedistributor_record5_payload_address;
assign main_rtio_core_outputs_record5_payload_data0 = main_rtio_core_outputs_lanedistributor_record5_payload_data;
assign main_rtio_core_outputs_record6_we = main_rtio_core_outputs_lanedistributor_record6_we;
assign main_rtio_core_outputs_lanedistributor_record6_writable = main_rtio_core_outputs_record6_writable;
assign main_rtio_core_outputs_record6_seqn0 = main_rtio_core_outputs_lanedistributor_record6_seqn;
assign main_rtio_core_outputs_record6_payload_channel0 = main_rtio_core_outputs_lanedistributor_record6_payload_channel;
assign main_rtio_core_outputs_record6_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
assign main_rtio_core_outputs_record6_payload_address0 = main_rtio_core_outputs_lanedistributor_record6_payload_address;
assign main_rtio_core_outputs_record6_payload_data0 = main_rtio_core_outputs_lanedistributor_record6_payload_data;
assign main_rtio_core_outputs_record7_we = main_rtio_core_outputs_lanedistributor_record7_we;
assign main_rtio_core_outputs_lanedistributor_record7_writable = main_rtio_core_outputs_record7_writable;
assign main_rtio_core_outputs_record7_seqn0 = main_rtio_core_outputs_lanedistributor_record7_seqn;
assign main_rtio_core_outputs_record7_payload_channel0 = main_rtio_core_outputs_lanedistributor_record7_payload_channel;
assign main_rtio_core_outputs_record7_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
assign main_rtio_core_outputs_record7_payload_address0 = main_rtio_core_outputs_lanedistributor_record7_payload_address;
assign main_rtio_core_outputs_record7_payload_data0 = main_rtio_core_outputs_lanedistributor_record7_payload_data;
assign main_rtio_core_outputs_record0_re = main_rtio_core_outputs_gates_record0_re;
assign main_rtio_core_outputs_gates_record0_readable = main_rtio_core_outputs_record0_readable;
assign main_rtio_core_outputs_gates_record0_seqn0 = main_rtio_core_outputs_record0_seqn1;
assign main_rtio_core_outputs_gates_record0_payload_channel0 = main_rtio_core_outputs_record0_payload_channel1;
assign main_rtio_core_outputs_gates_record0_payload_timestamp = main_rtio_core_outputs_record0_payload_timestamp1;
assign main_rtio_core_outputs_gates_record0_payload_address0 = main_rtio_core_outputs_record0_payload_address1;
assign main_rtio_core_outputs_gates_record0_payload_data0 = main_rtio_core_outputs_record0_payload_data1;
assign main_rtio_core_outputs_record1_re = main_rtio_core_outputs_gates_record1_re;
assign main_rtio_core_outputs_gates_record1_readable = main_rtio_core_outputs_record1_readable;
assign main_rtio_core_outputs_gates_record1_seqn0 = main_rtio_core_outputs_record1_seqn1;
assign main_rtio_core_outputs_gates_record1_payload_channel0 = main_rtio_core_outputs_record1_payload_channel1;
assign main_rtio_core_outputs_gates_record1_payload_timestamp = main_rtio_core_outputs_record1_payload_timestamp1;
assign main_rtio_core_outputs_gates_record1_payload_address0 = main_rtio_core_outputs_record1_payload_address1;
assign main_rtio_core_outputs_gates_record1_payload_data0 = main_rtio_core_outputs_record1_payload_data1;
assign main_rtio_core_outputs_record2_re = main_rtio_core_outputs_gates_record2_re;
assign main_rtio_core_outputs_gates_record2_readable = main_rtio_core_outputs_record2_readable;
assign main_rtio_core_outputs_gates_record2_seqn0 = main_rtio_core_outputs_record2_seqn1;
assign main_rtio_core_outputs_gates_record2_payload_channel0 = main_rtio_core_outputs_record2_payload_channel1;
assign main_rtio_core_outputs_gates_record2_payload_timestamp = main_rtio_core_outputs_record2_payload_timestamp1;
assign main_rtio_core_outputs_gates_record2_payload_address0 = main_rtio_core_outputs_record2_payload_address1;
assign main_rtio_core_outputs_gates_record2_payload_data0 = main_rtio_core_outputs_record2_payload_data1;
assign main_rtio_core_outputs_record3_re = main_rtio_core_outputs_gates_record3_re;
assign main_rtio_core_outputs_gates_record3_readable = main_rtio_core_outputs_record3_readable;
assign main_rtio_core_outputs_gates_record3_seqn0 = main_rtio_core_outputs_record3_seqn1;
assign main_rtio_core_outputs_gates_record3_payload_channel0 = main_rtio_core_outputs_record3_payload_channel1;
assign main_rtio_core_outputs_gates_record3_payload_timestamp = main_rtio_core_outputs_record3_payload_timestamp1;
assign main_rtio_core_outputs_gates_record3_payload_address0 = main_rtio_core_outputs_record3_payload_address1;
assign main_rtio_core_outputs_gates_record3_payload_data0 = main_rtio_core_outputs_record3_payload_data1;
assign main_rtio_core_outputs_record4_re = main_rtio_core_outputs_gates_record4_re;
assign main_rtio_core_outputs_gates_record4_readable = main_rtio_core_outputs_record4_readable;
assign main_rtio_core_outputs_gates_record4_seqn0 = main_rtio_core_outputs_record4_seqn1;
assign main_rtio_core_outputs_gates_record4_payload_channel0 = main_rtio_core_outputs_record4_payload_channel1;
assign main_rtio_core_outputs_gates_record4_payload_timestamp = main_rtio_core_outputs_record4_payload_timestamp1;
assign main_rtio_core_outputs_gates_record4_payload_address0 = main_rtio_core_outputs_record4_payload_address1;
assign main_rtio_core_outputs_gates_record4_payload_data0 = main_rtio_core_outputs_record4_payload_data1;
assign main_rtio_core_outputs_record5_re = main_rtio_core_outputs_gates_record5_re;
assign main_rtio_core_outputs_gates_record5_readable = main_rtio_core_outputs_record5_readable;
assign main_rtio_core_outputs_gates_record5_seqn0 = main_rtio_core_outputs_record5_seqn1;
assign main_rtio_core_outputs_gates_record5_payload_channel0 = main_rtio_core_outputs_record5_payload_channel1;
assign main_rtio_core_outputs_gates_record5_payload_timestamp = main_rtio_core_outputs_record5_payload_timestamp1;
assign main_rtio_core_outputs_gates_record5_payload_address0 = main_rtio_core_outputs_record5_payload_address1;
assign main_rtio_core_outputs_gates_record5_payload_data0 = main_rtio_core_outputs_record5_payload_data1;
assign main_rtio_core_outputs_record6_re = main_rtio_core_outputs_gates_record6_re;
assign main_rtio_core_outputs_gates_record6_readable = main_rtio_core_outputs_record6_readable;
assign main_rtio_core_outputs_gates_record6_seqn0 = main_rtio_core_outputs_record6_seqn1;
assign main_rtio_core_outputs_gates_record6_payload_channel0 = main_rtio_core_outputs_record6_payload_channel1;
assign main_rtio_core_outputs_gates_record6_payload_timestamp = main_rtio_core_outputs_record6_payload_timestamp1;
assign main_rtio_core_outputs_gates_record6_payload_address0 = main_rtio_core_outputs_record6_payload_address1;
assign main_rtio_core_outputs_gates_record6_payload_data0 = main_rtio_core_outputs_record6_payload_data1;
assign main_rtio_core_outputs_record7_re = main_rtio_core_outputs_gates_record7_re;
assign main_rtio_core_outputs_gates_record7_readable = main_rtio_core_outputs_record7_readable;
assign main_rtio_core_outputs_gates_record7_seqn0 = main_rtio_core_outputs_record7_seqn1;
assign main_rtio_core_outputs_gates_record7_payload_channel0 = main_rtio_core_outputs_record7_payload_channel1;
assign main_rtio_core_outputs_gates_record7_payload_timestamp = main_rtio_core_outputs_record7_payload_timestamp1;
assign main_rtio_core_outputs_gates_record7_payload_address0 = main_rtio_core_outputs_record7_payload_address1;
assign main_rtio_core_outputs_gates_record7_payload_data0 = main_rtio_core_outputs_record7_payload_data1;
assign main_rtio_core_outputs_record0_valid0 = main_rtio_core_outputs_gates_record0_valid;
assign main_rtio_core_outputs_record0_seqn2 = main_rtio_core_outputs_gates_record0_seqn1;
assign main_rtio_core_outputs_record0_replace_occured = main_rtio_core_outputs_gates_record0_replace_occured;
assign main_rtio_core_outputs_record0_nondata_replace_occured = main_rtio_core_outputs_gates_record0_nondata_replace_occured;
assign main_rtio_core_outputs_record0_payload_channel2 = main_rtio_core_outputs_gates_record0_payload_channel1;
assign main_rtio_core_outputs_record0_payload_fine_ts0 = main_rtio_core_outputs_gates_record0_payload_fine_ts;
assign main_rtio_core_outputs_record0_payload_address2 = main_rtio_core_outputs_gates_record0_payload_address1;
assign main_rtio_core_outputs_record0_payload_data2 = main_rtio_core_outputs_gates_record0_payload_data1;
assign main_rtio_core_outputs_record1_valid0 = main_rtio_core_outputs_gates_record1_valid;
assign main_rtio_core_outputs_record1_seqn2 = main_rtio_core_outputs_gates_record1_seqn1;
assign main_rtio_core_outputs_record1_replace_occured = main_rtio_core_outputs_gates_record1_replace_occured;
assign main_rtio_core_outputs_record1_nondata_replace_occured = main_rtio_core_outputs_gates_record1_nondata_replace_occured;
assign main_rtio_core_outputs_record1_payload_channel2 = main_rtio_core_outputs_gates_record1_payload_channel1;
assign main_rtio_core_outputs_record1_payload_fine_ts0 = main_rtio_core_outputs_gates_record1_payload_fine_ts;
assign main_rtio_core_outputs_record1_payload_address2 = main_rtio_core_outputs_gates_record1_payload_address1;
assign main_rtio_core_outputs_record1_payload_data2 = main_rtio_core_outputs_gates_record1_payload_data1;
assign main_rtio_core_outputs_record2_valid0 = main_rtio_core_outputs_gates_record2_valid;
assign main_rtio_core_outputs_record2_seqn2 = main_rtio_core_outputs_gates_record2_seqn1;
assign main_rtio_core_outputs_record2_replace_occured = main_rtio_core_outputs_gates_record2_replace_occured;
assign main_rtio_core_outputs_record2_nondata_replace_occured = main_rtio_core_outputs_gates_record2_nondata_replace_occured;
assign main_rtio_core_outputs_record2_payload_channel2 = main_rtio_core_outputs_gates_record2_payload_channel1;
assign main_rtio_core_outputs_record2_payload_fine_ts0 = main_rtio_core_outputs_gates_record2_payload_fine_ts;
assign main_rtio_core_outputs_record2_payload_address2 = main_rtio_core_outputs_gates_record2_payload_address1;
assign main_rtio_core_outputs_record2_payload_data2 = main_rtio_core_outputs_gates_record2_payload_data1;
assign main_rtio_core_outputs_record3_valid0 = main_rtio_core_outputs_gates_record3_valid;
assign main_rtio_core_outputs_record3_seqn2 = main_rtio_core_outputs_gates_record3_seqn1;
assign main_rtio_core_outputs_record3_replace_occured = main_rtio_core_outputs_gates_record3_replace_occured;
assign main_rtio_core_outputs_record3_nondata_replace_occured = main_rtio_core_outputs_gates_record3_nondata_replace_occured;
assign main_rtio_core_outputs_record3_payload_channel2 = main_rtio_core_outputs_gates_record3_payload_channel1;
assign main_rtio_core_outputs_record3_payload_fine_ts0 = main_rtio_core_outputs_gates_record3_payload_fine_ts;
assign main_rtio_core_outputs_record3_payload_address2 = main_rtio_core_outputs_gates_record3_payload_address1;
assign main_rtio_core_outputs_record3_payload_data2 = main_rtio_core_outputs_gates_record3_payload_data1;
assign main_rtio_core_outputs_record4_valid0 = main_rtio_core_outputs_gates_record4_valid;
assign main_rtio_core_outputs_record4_seqn2 = main_rtio_core_outputs_gates_record4_seqn1;
assign main_rtio_core_outputs_record4_replace_occured = main_rtio_core_outputs_gates_record4_replace_occured;
assign main_rtio_core_outputs_record4_nondata_replace_occured = main_rtio_core_outputs_gates_record4_nondata_replace_occured;
assign main_rtio_core_outputs_record4_payload_channel2 = main_rtio_core_outputs_gates_record4_payload_channel1;
assign main_rtio_core_outputs_record4_payload_fine_ts0 = main_rtio_core_outputs_gates_record4_payload_fine_ts;
assign main_rtio_core_outputs_record4_payload_address2 = main_rtio_core_outputs_gates_record4_payload_address1;
assign main_rtio_core_outputs_record4_payload_data2 = main_rtio_core_outputs_gates_record4_payload_data1;
assign main_rtio_core_outputs_record5_valid0 = main_rtio_core_outputs_gates_record5_valid;
assign main_rtio_core_outputs_record5_seqn2 = main_rtio_core_outputs_gates_record5_seqn1;
assign main_rtio_core_outputs_record5_replace_occured = main_rtio_core_outputs_gates_record5_replace_occured;
assign main_rtio_core_outputs_record5_nondata_replace_occured = main_rtio_core_outputs_gates_record5_nondata_replace_occured;
assign main_rtio_core_outputs_record5_payload_channel2 = main_rtio_core_outputs_gates_record5_payload_channel1;
assign main_rtio_core_outputs_record5_payload_fine_ts0 = main_rtio_core_outputs_gates_record5_payload_fine_ts;
assign main_rtio_core_outputs_record5_payload_address2 = main_rtio_core_outputs_gates_record5_payload_address1;
assign main_rtio_core_outputs_record5_payload_data2 = main_rtio_core_outputs_gates_record5_payload_data1;
assign main_rtio_core_outputs_record6_valid0 = main_rtio_core_outputs_gates_record6_valid;
assign main_rtio_core_outputs_record6_seqn2 = main_rtio_core_outputs_gates_record6_seqn1;
assign main_rtio_core_outputs_record6_replace_occured = main_rtio_core_outputs_gates_record6_replace_occured;
assign main_rtio_core_outputs_record6_nondata_replace_occured = main_rtio_core_outputs_gates_record6_nondata_replace_occured;
assign main_rtio_core_outputs_record6_payload_channel2 = main_rtio_core_outputs_gates_record6_payload_channel1;
assign main_rtio_core_outputs_record6_payload_fine_ts0 = main_rtio_core_outputs_gates_record6_payload_fine_ts;
assign main_rtio_core_outputs_record6_payload_address2 = main_rtio_core_outputs_gates_record6_payload_address1;
assign main_rtio_core_outputs_record6_payload_data2 = main_rtio_core_outputs_gates_record6_payload_data1;
assign main_rtio_core_outputs_record7_valid0 = main_rtio_core_outputs_gates_record7_valid;
assign main_rtio_core_outputs_record7_seqn2 = main_rtio_core_outputs_gates_record7_seqn1;
assign main_rtio_core_outputs_record7_replace_occured = main_rtio_core_outputs_gates_record7_replace_occured;
assign main_rtio_core_outputs_record7_nondata_replace_occured = main_rtio_core_outputs_gates_record7_nondata_replace_occured;
assign main_rtio_core_outputs_record7_payload_channel2 = main_rtio_core_outputs_gates_record7_payload_channel1;
assign main_rtio_core_outputs_record7_payload_fine_ts0 = main_rtio_core_outputs_gates_record7_payload_fine_ts;
assign main_rtio_core_outputs_record7_payload_address2 = main_rtio_core_outputs_gates_record7_payload_address1;
assign main_rtio_core_outputs_record7_payload_data2 = main_rtio_core_outputs_gates_record7_payload_data1;
assign main_rtio_core_cri_o_status = {main_rtio_core_outputs_lanedistributor_o_status_underflow, main_rtio_core_outputs_lanedistributor_o_status_wait};
assign main_rtio_core_outputs_lanedistributor_record0_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record0_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record0_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record0_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record1_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record1_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record1_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record1_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record2_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record2_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record2_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record2_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record3_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record3_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record3_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record3_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record4_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record4_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record4_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record4_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record5_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record5_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record5_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record5_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record6_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record6_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record6_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record6_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record7_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record7_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record7_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record7_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_coarse_timestamp = main_rtio_core_cri_o_timestamp[63:3];
assign main_rtio_core_outputs_lanedistributor_current_lane_plus_one = (main_rtio_core_outputs_lanedistributor_current_lane + 1'd1);
assign main_rtio_core_outputs_lanedistributor_adr = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_compensation = main_rtio_core_outputs_lanedistributor_dat_r;
assign main_rtio_core_outputs_lanedistributor_timestamp_above_min = ((main_rtio_core_outputs_lanedistributor_min_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min = ((main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min = ((main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_last = ((main_rtio_core_outputs_lanedistributor_last_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));

// synthesis translate_off
reg dummy_d_86;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	main_rtio_core_outputs_lanedistributor_use_lanen <= 3'd0;
	if ((main_rtio_core_outputs_lanedistributor_force_laneB | (~main_rtio_core_outputs_lanedistributor_timestamp_above_last))) begin
		main_rtio_core_outputs_lanedistributor_use_lanen <= main_rtio_core_outputs_lanedistributor_current_lane_plus_one;
		main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd1;
	end else begin
		main_rtio_core_outputs_lanedistributor_use_lanen <= main_rtio_core_outputs_lanedistributor_current_lane;
		main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	end
// synthesis translate_off
	dummy_d_86 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min = (main_rtio_core_outputs_lanedistributor_use_laneB ? main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min : main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min);

// synthesis translate_off
reg dummy_d_87;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_do_write <= 1'd0;
	main_rtio_core_outputs_lanedistributor_do_underflow <= 1'd0;
	main_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd0;
	if (((~main_rtio_core_outputs_lanedistributor_quash) & (main_rtio_core_cri_cmd == 1'd1))) begin
		if (main_rtio_core_outputs_lanedistributor_timestamp_above_min) begin
			if (main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min) begin
				main_rtio_core_outputs_lanedistributor_do_write <= 1'd1;
			end else begin
				main_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd1;
			end
		end else begin
			main_rtio_core_outputs_lanedistributor_do_underflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_87 <= dummy_s;
// synthesis translate_on
end
assign builder_comb_lhs_array_muxed = main_rtio_core_outputs_lanedistributor_do_write;

// synthesis translate_off
reg dummy_d_88;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record0_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record1_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record2_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record3_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record4_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record5_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record6_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record7_we <= 1'd0;
	case (main_rtio_core_outputs_lanedistributor_use_lanen)
		1'd0: begin
			main_rtio_core_outputs_lanedistributor_record0_we <= builder_comb_lhs_array_muxed;
		end
		1'd1: begin
			main_rtio_core_outputs_lanedistributor_record1_we <= builder_comb_lhs_array_muxed;
		end
		2'd2: begin
			main_rtio_core_outputs_lanedistributor_record2_we <= builder_comb_lhs_array_muxed;
		end
		2'd3: begin
			main_rtio_core_outputs_lanedistributor_record3_we <= builder_comb_lhs_array_muxed;
		end
		3'd4: begin
			main_rtio_core_outputs_lanedistributor_record4_we <= builder_comb_lhs_array_muxed;
		end
		3'd5: begin
			main_rtio_core_outputs_lanedistributor_record5_we <= builder_comb_lhs_array_muxed;
		end
		3'd6: begin
			main_rtio_core_outputs_lanedistributor_record6_we <= builder_comb_lhs_array_muxed;
		end
		default: begin
			main_rtio_core_outputs_lanedistributor_record7_we <= builder_comb_lhs_array_muxed;
		end
	endcase
// synthesis translate_off
	dummy_d_88 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_compensated_timestamp = ($signed({1'd0, main_rtio_core_cri_o_timestamp}) + (main_rtio_core_outputs_lanedistributor_compensation <<< 2'd3));

// synthesis translate_off
reg dummy_d_89;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_89 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_90;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_90 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_91;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_91 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_92;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_92 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_93;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_93 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_94;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_94 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_95;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_95 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_96;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_96 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_current_lane_writable = builder_comb_rhs_array_muxed8;
assign main_rtio_core_outputs_lanedistributor_o_status_wait = (~main_rtio_core_outputs_lanedistributor_current_lane_writable);
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din = {{main_rtio_core_outputs_record0_payload_data0, main_rtio_core_outputs_record0_payload_address0, main_rtio_core_outputs_record0_payload_timestamp0, main_rtio_core_outputs_record0_payload_channel0}, main_rtio_core_outputs_record0_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we = main_rtio_core_outputs_record0_we;
assign main_rtio_core_outputs_record0_writable = main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
assign {{main_rtio_core_outputs_record0_payload_data1, main_rtio_core_outputs_record0_payload_address1, main_rtio_core_outputs_record0_payload_timestamp1, main_rtio_core_outputs_record0_payload_channel1}, main_rtio_core_outputs_record0_seqn1} = main_rtio_core_outputs_asyncfifobuffered0_dout;
assign main_rtio_core_outputs_record0_readable = main_rtio_core_outputs_asyncfifobuffered0_readable;
assign main_rtio_core_outputs_asyncfifobuffered0_re = main_rtio_core_outputs_record0_re;
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din = {{main_rtio_core_outputs_record1_payload_data0, main_rtio_core_outputs_record1_payload_address0, main_rtio_core_outputs_record1_payload_timestamp0, main_rtio_core_outputs_record1_payload_channel0}, main_rtio_core_outputs_record1_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we = main_rtio_core_outputs_record1_we;
assign main_rtio_core_outputs_record1_writable = main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
assign {{main_rtio_core_outputs_record1_payload_data1, main_rtio_core_outputs_record1_payload_address1, main_rtio_core_outputs_record1_payload_timestamp1, main_rtio_core_outputs_record1_payload_channel1}, main_rtio_core_outputs_record1_seqn1} = main_rtio_core_outputs_asyncfifobuffered1_dout;
assign main_rtio_core_outputs_record1_readable = main_rtio_core_outputs_asyncfifobuffered1_readable;
assign main_rtio_core_outputs_asyncfifobuffered1_re = main_rtio_core_outputs_record1_re;
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din = {{main_rtio_core_outputs_record2_payload_data0, main_rtio_core_outputs_record2_payload_address0, main_rtio_core_outputs_record2_payload_timestamp0, main_rtio_core_outputs_record2_payload_channel0}, main_rtio_core_outputs_record2_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we = main_rtio_core_outputs_record2_we;
assign main_rtio_core_outputs_record2_writable = main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
assign {{main_rtio_core_outputs_record2_payload_data1, main_rtio_core_outputs_record2_payload_address1, main_rtio_core_outputs_record2_payload_timestamp1, main_rtio_core_outputs_record2_payload_channel1}, main_rtio_core_outputs_record2_seqn1} = main_rtio_core_outputs_asyncfifobuffered2_dout;
assign main_rtio_core_outputs_record2_readable = main_rtio_core_outputs_asyncfifobuffered2_readable;
assign main_rtio_core_outputs_asyncfifobuffered2_re = main_rtio_core_outputs_record2_re;
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din = {{main_rtio_core_outputs_record3_payload_data0, main_rtio_core_outputs_record3_payload_address0, main_rtio_core_outputs_record3_payload_timestamp0, main_rtio_core_outputs_record3_payload_channel0}, main_rtio_core_outputs_record3_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we = main_rtio_core_outputs_record3_we;
assign main_rtio_core_outputs_record3_writable = main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
assign {{main_rtio_core_outputs_record3_payload_data1, main_rtio_core_outputs_record3_payload_address1, main_rtio_core_outputs_record3_payload_timestamp1, main_rtio_core_outputs_record3_payload_channel1}, main_rtio_core_outputs_record3_seqn1} = main_rtio_core_outputs_asyncfifobuffered3_dout;
assign main_rtio_core_outputs_record3_readable = main_rtio_core_outputs_asyncfifobuffered3_readable;
assign main_rtio_core_outputs_asyncfifobuffered3_re = main_rtio_core_outputs_record3_re;
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din = {{main_rtio_core_outputs_record4_payload_data0, main_rtio_core_outputs_record4_payload_address0, main_rtio_core_outputs_record4_payload_timestamp0, main_rtio_core_outputs_record4_payload_channel0}, main_rtio_core_outputs_record4_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we = main_rtio_core_outputs_record4_we;
assign main_rtio_core_outputs_record4_writable = main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
assign {{main_rtio_core_outputs_record4_payload_data1, main_rtio_core_outputs_record4_payload_address1, main_rtio_core_outputs_record4_payload_timestamp1, main_rtio_core_outputs_record4_payload_channel1}, main_rtio_core_outputs_record4_seqn1} = main_rtio_core_outputs_asyncfifobuffered4_dout;
assign main_rtio_core_outputs_record4_readable = main_rtio_core_outputs_asyncfifobuffered4_readable;
assign main_rtio_core_outputs_asyncfifobuffered4_re = main_rtio_core_outputs_record4_re;
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din = {{main_rtio_core_outputs_record5_payload_data0, main_rtio_core_outputs_record5_payload_address0, main_rtio_core_outputs_record5_payload_timestamp0, main_rtio_core_outputs_record5_payload_channel0}, main_rtio_core_outputs_record5_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we = main_rtio_core_outputs_record5_we;
assign main_rtio_core_outputs_record5_writable = main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
assign {{main_rtio_core_outputs_record5_payload_data1, main_rtio_core_outputs_record5_payload_address1, main_rtio_core_outputs_record5_payload_timestamp1, main_rtio_core_outputs_record5_payload_channel1}, main_rtio_core_outputs_record5_seqn1} = main_rtio_core_outputs_asyncfifobuffered5_dout;
assign main_rtio_core_outputs_record5_readable = main_rtio_core_outputs_asyncfifobuffered5_readable;
assign main_rtio_core_outputs_asyncfifobuffered5_re = main_rtio_core_outputs_record5_re;
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din = {{main_rtio_core_outputs_record6_payload_data0, main_rtio_core_outputs_record6_payload_address0, main_rtio_core_outputs_record6_payload_timestamp0, main_rtio_core_outputs_record6_payload_channel0}, main_rtio_core_outputs_record6_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we = main_rtio_core_outputs_record6_we;
assign main_rtio_core_outputs_record6_writable = main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
assign {{main_rtio_core_outputs_record6_payload_data1, main_rtio_core_outputs_record6_payload_address1, main_rtio_core_outputs_record6_payload_timestamp1, main_rtio_core_outputs_record6_payload_channel1}, main_rtio_core_outputs_record6_seqn1} = main_rtio_core_outputs_asyncfifobuffered6_dout;
assign main_rtio_core_outputs_record6_readable = main_rtio_core_outputs_asyncfifobuffered6_readable;
assign main_rtio_core_outputs_asyncfifobuffered6_re = main_rtio_core_outputs_record6_re;
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din = {{main_rtio_core_outputs_record7_payload_data0, main_rtio_core_outputs_record7_payload_address0, main_rtio_core_outputs_record7_payload_timestamp0, main_rtio_core_outputs_record7_payload_channel0}, main_rtio_core_outputs_record7_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we = main_rtio_core_outputs_record7_we;
assign main_rtio_core_outputs_record7_writable = main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
assign {{main_rtio_core_outputs_record7_payload_data1, main_rtio_core_outputs_record7_payload_address1, main_rtio_core_outputs_record7_payload_timestamp1, main_rtio_core_outputs_record7_payload_channel1}, main_rtio_core_outputs_record7_seqn1} = main_rtio_core_outputs_asyncfifobuffered7_dout;
assign main_rtio_core_outputs_record7_readable = main_rtio_core_outputs_asyncfifobuffered7_readable;
assign main_rtio_core_outputs_asyncfifobuffered7_re = main_rtio_core_outputs_record7_re;
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re = (main_rtio_core_outputs_asyncfifobuffered0_re | (~main_rtio_core_outputs_asyncfifobuffered0_readable));
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce = (main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable & main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we);
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce = (main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable & main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re);
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable = (((main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[7] == main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[6] == main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[5:0] != main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable = (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q != main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_adr = main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_we = main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
assign main_rtio_core_outputs_asyncfifobuffered0_rdport_adr = main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout = main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_97;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce) begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_97 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next = (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_98;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce) begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_98 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next = (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re = (main_rtio_core_outputs_asyncfifobuffered1_re | (~main_rtio_core_outputs_asyncfifobuffered1_readable));
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce = (main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable & main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we);
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce = (main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable & main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re);
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable = (((main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[7] == main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[6] == main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[5:0] != main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable = (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q != main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_adr = main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_we = main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
assign main_rtio_core_outputs_asyncfifobuffered1_rdport_adr = main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout = main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_99;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce) begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_99 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next = (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_100;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce) begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_100 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next = (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re = (main_rtio_core_outputs_asyncfifobuffered2_re | (~main_rtio_core_outputs_asyncfifobuffered2_readable));
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce = (main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable & main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we);
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce = (main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable & main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re);
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable = (((main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[7] == main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[6] == main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[5:0] != main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable = (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q != main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_adr = main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_we = main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
assign main_rtio_core_outputs_asyncfifobuffered2_rdport_adr = main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout = main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_101;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce) begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_101 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next = (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_102;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce) begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_102 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next = (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re = (main_rtio_core_outputs_asyncfifobuffered3_re | (~main_rtio_core_outputs_asyncfifobuffered3_readable));
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce = (main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable & main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we);
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce = (main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable & main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re);
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable = (((main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[7] == main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[6] == main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[5:0] != main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable = (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q != main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_adr = main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_we = main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
assign main_rtio_core_outputs_asyncfifobuffered3_rdport_adr = main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout = main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_103;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce) begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_103 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next = (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_104;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce) begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_104 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next = (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re = (main_rtio_core_outputs_asyncfifobuffered4_re | (~main_rtio_core_outputs_asyncfifobuffered4_readable));
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce = (main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable & main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we);
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce = (main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable & main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re);
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable = (((main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[7] == main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[6] == main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[5:0] != main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable = (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q != main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_adr = main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_we = main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
assign main_rtio_core_outputs_asyncfifobuffered4_rdport_adr = main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout = main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_105;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce) begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_105 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next = (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_106;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce) begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_106 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next = (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re = (main_rtio_core_outputs_asyncfifobuffered5_re | (~main_rtio_core_outputs_asyncfifobuffered5_readable));
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce = (main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable & main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we);
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce = (main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable & main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re);
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable = (((main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[7] == main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[6] == main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[5:0] != main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable = (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q != main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_adr = main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_we = main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
assign main_rtio_core_outputs_asyncfifobuffered5_rdport_adr = main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout = main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_107;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce) begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_107 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next = (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_108;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce) begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_108 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next = (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re = (main_rtio_core_outputs_asyncfifobuffered6_re | (~main_rtio_core_outputs_asyncfifobuffered6_readable));
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce = (main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable & main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we);
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce = (main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable & main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re);
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable = (((main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[7] == main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[6] == main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[5:0] != main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable = (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q != main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_adr = main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_we = main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
assign main_rtio_core_outputs_asyncfifobuffered6_rdport_adr = main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout = main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_109;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce) begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_109 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next = (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_110;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce) begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_110 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next = (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re = (main_rtio_core_outputs_asyncfifobuffered7_re | (~main_rtio_core_outputs_asyncfifobuffered7_readable));
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce = (main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable & main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we);
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce = (main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable & main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re);
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable = (((main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[7] == main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[6] == main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[5:0] != main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable = (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q != main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_adr = main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_we = main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
assign main_rtio_core_outputs_asyncfifobuffered7_rdport_adr = main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout = main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;

// synthesis translate_off
reg dummy_d_111;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce) begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary;
	end
// synthesis translate_off
	dummy_d_111 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next = (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_112;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce) begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary;
	end
// synthesis translate_off
	dummy_d_112 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next = (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[7:1]);
assign main_rtio_core_outputs_gates_record0_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record0_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record0_re = (main_rtio_core_outputs_gates_record0_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record1_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record1_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record1_re = (main_rtio_core_outputs_gates_record1_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record2_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record2_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record2_re = (main_rtio_core_outputs_gates_record2_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record3_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record3_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record3_re = (main_rtio_core_outputs_gates_record3_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record4_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record4_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record4_re = (main_rtio_core_outputs_gates_record4_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record5_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record5_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record5_re = (main_rtio_core_outputs_gates_record5_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record6_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record6_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record6_re = (main_rtio_core_outputs_gates_record6_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record7_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record7_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record7_re = (main_rtio_core_outputs_gates_record7_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_memory0_adr = main_rtio_core_outputs_record40_rec_payload_channel;
assign main_rtio_core_outputs_record0_collision = (main_rtio_core_outputs_replace_occured_r0 & ((~main_rtio_core_outputs_memory0_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r0));
assign main_rtio_core_outputs_memory1_adr = main_rtio_core_outputs_record41_rec_payload_channel;
assign main_rtio_core_outputs_record1_collision = (main_rtio_core_outputs_replace_occured_r1 & ((~main_rtio_core_outputs_memory1_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r1));
assign main_rtio_core_outputs_memory2_adr = main_rtio_core_outputs_record42_rec_payload_channel;
assign main_rtio_core_outputs_record2_collision = (main_rtio_core_outputs_replace_occured_r2 & ((~main_rtio_core_outputs_memory2_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r2));
assign main_rtio_core_outputs_memory3_adr = main_rtio_core_outputs_record43_rec_payload_channel;
assign main_rtio_core_outputs_record3_collision = (main_rtio_core_outputs_replace_occured_r3 & ((~main_rtio_core_outputs_memory3_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r3));
assign main_rtio_core_outputs_memory4_adr = main_rtio_core_outputs_record44_rec_payload_channel;
assign main_rtio_core_outputs_record4_collision = (main_rtio_core_outputs_replace_occured_r4 & ((~main_rtio_core_outputs_memory4_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r4));
assign main_rtio_core_outputs_memory5_adr = main_rtio_core_outputs_record45_rec_payload_channel;
assign main_rtio_core_outputs_record5_collision = (main_rtio_core_outputs_replace_occured_r5 & ((~main_rtio_core_outputs_memory5_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r5));
assign main_rtio_core_outputs_memory6_adr = main_rtio_core_outputs_record46_rec_payload_channel;
assign main_rtio_core_outputs_record6_collision = (main_rtio_core_outputs_replace_occured_r6 & ((~main_rtio_core_outputs_memory6_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r6));
assign main_rtio_core_outputs_memory7_adr = main_rtio_core_outputs_record47_rec_payload_channel;
assign main_rtio_core_outputs_record7_collision = (main_rtio_core_outputs_replace_occured_r7 & ((~main_rtio_core_outputs_memory7_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r7));
assign main_rtio_core_outputs_selected0 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected1 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected2 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected3 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected4 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected5 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected6 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected7 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected8 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected9 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected10 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected11 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected12 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected13 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected14 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected15 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected16 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected17 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected18 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected19 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected20 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected21 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected22 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected23 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected24 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected25 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected26 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected27 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected28 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected29 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected30 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected31 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected32 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected33 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected34 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected35 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected36 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected37 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected38 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected39 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected40 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected41 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected42 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected43 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected44 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected45 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected46 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected47 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected48 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected49 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected50 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected51 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected52 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected53 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected54 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected55 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected56 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected57 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected58 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected59 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected60 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected61 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected62 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected63 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected64 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected65 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected66 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected67 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected68 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected69 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected70 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected71 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected72 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected73 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected74 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected75 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected76 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected77 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected78 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected79 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected80 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected81 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected82 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected83 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected84 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected85 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected86 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected87 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected88 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected89 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected90 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected91 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected92 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected93 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected94 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected95 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected96 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected97 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected98 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected99 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected100 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected101 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected102 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected103 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected104 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected105 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected106 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected107 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected108 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected109 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected110 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected111 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected112 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected113 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected114 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected115 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected116 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected117 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected118 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected119 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected120 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected121 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected122 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected123 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected124 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected125 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected126 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected127 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected128 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected129 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected130 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected131 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected132 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected133 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected134 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected135 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected136 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected137 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected138 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected139 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected140 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected141 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected142 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected143 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected144 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected145 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected146 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected147 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected148 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected149 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected150 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected151 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected152 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected153 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected154 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected155 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected156 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected157 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected158 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected159 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected160 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected161 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected162 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected163 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected164 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected165 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected166 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected167 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected168 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected169 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected170 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected171 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected172 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected173 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected174 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected175 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected176 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected177 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected178 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected179 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected180 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected181 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected182 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected183 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected184 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected185 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected186 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected187 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected188 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected189 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected190 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected191 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected192 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected193 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected194 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected195 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected196 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected197 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected198 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected199 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected200 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected201 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected202 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected203 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected204 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected205 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected206 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected207 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected208 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected209 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected210 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected211 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected212 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected213 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected214 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected215 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected216 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected217 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected218 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected219 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected220 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected221 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected222 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected223 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected224 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected225 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected226 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected227 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected228 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected229 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected230 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected231 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected232 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected233 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected234 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected235 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected236 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected237 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected238 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected239 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd29));
assign main_rtio_core_outputs_selected240 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected241 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected242 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected243 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected244 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected245 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected246 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected247 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd30));
assign main_rtio_core_outputs_selected248 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected249 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected250 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected251 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected252 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected253 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected254 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected255 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd31));
assign main_rtio_core_outputs_selected256 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected257 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected258 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected259 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected260 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected261 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected262 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected263 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 6'd32));
assign main_rtio_core_outputs_selected264 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected265 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected266 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected267 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected268 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected269 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected270 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected271 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 6'd33));
assign main_rtio_core_outputs_selected272 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected273 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected274 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected275 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected276 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected277 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected278 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected279 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 6'd34));
assign main_rtio_core_outputs_selected280 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected281 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected282 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected283 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected284 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected285 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected286 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected287 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 6'd35));
assign main_rtio_core_outputs_selected288 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected289 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected290 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected291 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected292 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected293 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected294 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 6'd36));
assign main_rtio_core_outputs_selected295 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 6'd36));

// synthesis translate_off
reg dummy_d_113;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference0 <= 1'd0;
	if ((main_rtio_core_outputs_record0_payload_channel2 != main_rtio_core_outputs_record1_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_payload_fine_ts0 != main_rtio_core_outputs_record1_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_payload_address2 != main_rtio_core_outputs_record1_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_113 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_114;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference1 <= 1'd0;
	if ((main_rtio_core_outputs_record2_payload_channel2 != main_rtio_core_outputs_record3_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record2_payload_fine_ts0 != main_rtio_core_outputs_record3_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record2_payload_address2 != main_rtio_core_outputs_record3_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_114 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_115;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference2 <= 1'd0;
	if ((main_rtio_core_outputs_record4_payload_channel2 != main_rtio_core_outputs_record5_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_payload_fine_ts0 != main_rtio_core_outputs_record5_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_payload_address2 != main_rtio_core_outputs_record5_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_115 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_116;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference3 <= 1'd0;
	if ((main_rtio_core_outputs_record6_payload_channel2 != main_rtio_core_outputs_record7_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record6_payload_fine_ts0 != main_rtio_core_outputs_record7_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record6_payload_address2 != main_rtio_core_outputs_record7_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_116 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_117;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference4 <= 1'd0;
	if ((main_rtio_core_outputs_record0_rec_payload_channel != main_rtio_core_outputs_record2_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_rec_payload_fine_ts != main_rtio_core_outputs_record2_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_rec_payload_address != main_rtio_core_outputs_record2_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_117 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_118;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference5 <= 1'd0;
	if ((main_rtio_core_outputs_record1_rec_payload_channel != main_rtio_core_outputs_record3_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record1_rec_payload_fine_ts != main_rtio_core_outputs_record3_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record1_rec_payload_address != main_rtio_core_outputs_record3_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_118 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_119;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference6 <= 1'd0;
	if ((main_rtio_core_outputs_record4_rec_payload_channel != main_rtio_core_outputs_record6_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_rec_payload_fine_ts != main_rtio_core_outputs_record6_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_rec_payload_address != main_rtio_core_outputs_record6_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_119 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_120;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference7 <= 1'd0;
	if ((main_rtio_core_outputs_record5_rec_payload_channel != main_rtio_core_outputs_record7_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record5_rec_payload_fine_ts != main_rtio_core_outputs_record7_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record5_rec_payload_address != main_rtio_core_outputs_record7_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_120 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_121;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference8 <= 1'd0;
	if ((main_rtio_core_outputs_record9_rec_payload_channel != main_rtio_core_outputs_record10_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record9_rec_payload_fine_ts != main_rtio_core_outputs_record10_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record9_rec_payload_address != main_rtio_core_outputs_record10_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_121 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_122;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference9 <= 1'd0;
	if ((main_rtio_core_outputs_record13_rec_payload_channel != main_rtio_core_outputs_record14_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record13_rec_payload_fine_ts != main_rtio_core_outputs_record14_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record13_rec_payload_address != main_rtio_core_outputs_record14_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_122 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_123;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference10 <= 1'd0;
	if ((main_rtio_core_outputs_record16_rec_payload_channel != main_rtio_core_outputs_record20_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record16_rec_payload_fine_ts != main_rtio_core_outputs_record20_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record16_rec_payload_address != main_rtio_core_outputs_record20_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_123 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_124;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference11 <= 1'd0;
	if ((main_rtio_core_outputs_record17_rec_payload_channel != main_rtio_core_outputs_record21_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record17_rec_payload_fine_ts != main_rtio_core_outputs_record21_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record17_rec_payload_address != main_rtio_core_outputs_record21_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_124 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_125;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference12 <= 1'd0;
	if ((main_rtio_core_outputs_record18_rec_payload_channel != main_rtio_core_outputs_record22_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record18_rec_payload_fine_ts != main_rtio_core_outputs_record22_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record18_rec_payload_address != main_rtio_core_outputs_record22_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_125 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_126;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference13 <= 1'd0;
	if ((main_rtio_core_outputs_record19_rec_payload_channel != main_rtio_core_outputs_record23_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record19_rec_payload_fine_ts != main_rtio_core_outputs_record23_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record19_rec_payload_address != main_rtio_core_outputs_record23_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_126 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_127;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference14 <= 1'd0;
	if ((main_rtio_core_outputs_record26_rec_payload_channel != main_rtio_core_outputs_record28_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record26_rec_payload_fine_ts != main_rtio_core_outputs_record28_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record26_rec_payload_address != main_rtio_core_outputs_record28_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_127 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_128;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference15 <= 1'd0;
	if ((main_rtio_core_outputs_record27_rec_payload_channel != main_rtio_core_outputs_record29_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record27_rec_payload_fine_ts != main_rtio_core_outputs_record29_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record27_rec_payload_address != main_rtio_core_outputs_record29_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_128 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_129;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference16 <= 1'd0;
	if ((main_rtio_core_outputs_record33_rec_payload_channel != main_rtio_core_outputs_record34_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record33_rec_payload_fine_ts != main_rtio_core_outputs_record34_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record33_rec_payload_address != main_rtio_core_outputs_record34_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_129 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_130;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference17 <= 1'd0;
	if ((main_rtio_core_outputs_record35_rec_payload_channel != main_rtio_core_outputs_record36_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record35_rec_payload_fine_ts != main_rtio_core_outputs_record36_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record35_rec_payload_address != main_rtio_core_outputs_record36_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_130 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_131;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference18 <= 1'd0;
	if ((main_rtio_core_outputs_record37_rec_payload_channel != main_rtio_core_outputs_record38_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record37_rec_payload_fine_ts != main_rtio_core_outputs_record38_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record37_rec_payload_address != main_rtio_core_outputs_record38_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_131 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_din = {main_rtio_core_inputs_record0_fifo_in_timestamp, main_rtio_core_inputs_record0_fifo_in_data};
assign {main_rtio_core_inputs_record0_fifo_out_timestamp, main_rtio_core_inputs_record0_fifo_out_data} = main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
assign main_rtio_core_inputs_record0_fifo_in_data = main_inout_8x0_inout_8x0_iinterface0_data;
assign main_rtio_core_inputs_record0_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x0_inout_8x0_iinterface0_fine_ts};
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_we = main_inout_8x0_inout_8x0_iinterface0_stb;
assign main_rtio_core_inputs_overflow_io0 = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_we & (~main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable));
assign main_rtio_core_inputs_blindtransfer0_i = main_rtio_core_inputs_overflow_io0;
assign main_rtio_core_inputs_selected0 = (main_rtio_core_cri_chan_sel[15:0] == 1'd0);
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_re = ((main_rtio_core_inputs_selected0 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow0));
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_din = {main_rtio_core_inputs_record1_fifo_in_timestamp, main_rtio_core_inputs_record1_fifo_in_data};
assign {main_rtio_core_inputs_record1_fifo_out_timestamp, main_rtio_core_inputs_record1_fifo_out_data} = main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
assign main_rtio_core_inputs_record1_fifo_in_data = main_inout_8x1_inout_8x1_iinterface1_data;
assign main_rtio_core_inputs_record1_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x1_inout_8x1_iinterface1_fine_ts};
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_we = main_inout_8x1_inout_8x1_iinterface1_stb;
assign main_rtio_core_inputs_overflow_io1 = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_we & (~main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable));
assign main_rtio_core_inputs_blindtransfer1_i = main_rtio_core_inputs_overflow_io1;
assign main_rtio_core_inputs_selected1 = (main_rtio_core_cri_chan_sel[15:0] == 1'd1);
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_re = ((main_rtio_core_inputs_selected1 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow1));
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_din = {main_rtio_core_inputs_record2_fifo_in_timestamp, main_rtio_core_inputs_record2_fifo_in_data};
assign {main_rtio_core_inputs_record2_fifo_out_timestamp, main_rtio_core_inputs_record2_fifo_out_data} = main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
assign main_rtio_core_inputs_record2_fifo_in_data = main_inout_8x2_inout_8x2_iinterface2_data;
assign main_rtio_core_inputs_record2_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x2_inout_8x2_iinterface2_fine_ts};
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_we = main_inout_8x2_inout_8x2_iinterface2_stb;
assign main_rtio_core_inputs_overflow_io2 = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_we & (~main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable));
assign main_rtio_core_inputs_blindtransfer2_i = main_rtio_core_inputs_overflow_io2;
assign main_rtio_core_inputs_selected2 = (main_rtio_core_cri_chan_sel[15:0] == 2'd2);
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_re = ((main_rtio_core_inputs_selected2 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow2));
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_din = {main_rtio_core_inputs_record3_fifo_in_timestamp, main_rtio_core_inputs_record3_fifo_in_data};
assign {main_rtio_core_inputs_record3_fifo_out_timestamp, main_rtio_core_inputs_record3_fifo_out_data} = main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
assign main_rtio_core_inputs_record3_fifo_in_data = main_inout_8x3_inout_8x3_iinterface3_data;
assign main_rtio_core_inputs_record3_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x3_inout_8x3_iinterface3_fine_ts};
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_we = main_inout_8x3_inout_8x3_iinterface3_stb;
assign main_rtio_core_inputs_overflow_io3 = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_we & (~main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable));
assign main_rtio_core_inputs_blindtransfer3_i = main_rtio_core_inputs_overflow_io3;
assign main_rtio_core_inputs_selected3 = (main_rtio_core_cri_chan_sel[15:0] == 2'd3);
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_re = ((main_rtio_core_inputs_selected3 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow3));
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_din = {main_rtio_core_inputs_record4_fifo_in_timestamp, main_rtio_core_inputs_record4_fifo_in_data};
assign {main_rtio_core_inputs_record4_fifo_out_timestamp, main_rtio_core_inputs_record4_fifo_out_data} = main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
assign main_rtio_core_inputs_record4_fifo_in_data = main_inout_8x4_inout_8x4_iinterface4_data;
assign main_rtio_core_inputs_record4_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x4_inout_8x4_iinterface4_fine_ts};
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_we = main_inout_8x4_inout_8x4_iinterface4_stb;
assign main_rtio_core_inputs_overflow_io4 = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_we & (~main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable));
assign main_rtio_core_inputs_blindtransfer4_i = main_rtio_core_inputs_overflow_io4;
assign main_rtio_core_inputs_selected4 = (main_rtio_core_cri_chan_sel[15:0] == 3'd4);
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_re = ((main_rtio_core_inputs_selected4 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow4));
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_din = {main_rtio_core_inputs_record5_fifo_in_timestamp, main_rtio_core_inputs_record5_fifo_in_data};
assign {main_rtio_core_inputs_record5_fifo_out_timestamp, main_rtio_core_inputs_record5_fifo_out_data} = main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
assign main_rtio_core_inputs_record5_fifo_in_data = main_inout_8x5_inout_8x5_iinterface5_data;
assign main_rtio_core_inputs_record5_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x5_inout_8x5_iinterface5_fine_ts};
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_we = main_inout_8x5_inout_8x5_iinterface5_stb;
assign main_rtio_core_inputs_overflow_io5 = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_we & (~main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable));
assign main_rtio_core_inputs_blindtransfer5_i = main_rtio_core_inputs_overflow_io5;
assign main_rtio_core_inputs_selected5 = (main_rtio_core_cri_chan_sel[15:0] == 3'd5);
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_re = ((main_rtio_core_inputs_selected5 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow5));
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_din = {main_rtio_core_inputs_record6_fifo_in_timestamp, main_rtio_core_inputs_record6_fifo_in_data};
assign {main_rtio_core_inputs_record6_fifo_out_timestamp, main_rtio_core_inputs_record6_fifo_out_data} = main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
assign main_rtio_core_inputs_record6_fifo_in_data = main_inout_8x6_inout_8x6_iinterface6_data;
assign main_rtio_core_inputs_record6_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x6_inout_8x6_iinterface6_fine_ts};
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_we = main_inout_8x6_inout_8x6_iinterface6_stb;
assign main_rtio_core_inputs_overflow_io6 = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_we & (~main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable));
assign main_rtio_core_inputs_blindtransfer6_i = main_rtio_core_inputs_overflow_io6;
assign main_rtio_core_inputs_selected6 = (main_rtio_core_cri_chan_sel[15:0] == 3'd6);
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_re = ((main_rtio_core_inputs_selected6 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow6));
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_din = {main_rtio_core_inputs_record7_fifo_in_timestamp, main_rtio_core_inputs_record7_fifo_in_data};
assign {main_rtio_core_inputs_record7_fifo_out_timestamp, main_rtio_core_inputs_record7_fifo_out_data} = main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout;
assign main_rtio_core_inputs_record7_fifo_in_data = main_inout_8x7_inout_8x7_iinterface7_data;
assign main_rtio_core_inputs_record7_fifo_in_timestamp = {main_rtio_tsc_coarse_ts, main_inout_8x7_inout_8x7_iinterface7_fine_ts};
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_we = main_inout_8x7_inout_8x7_iinterface7_stb;
assign main_rtio_core_inputs_overflow_io7 = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_we & (~main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable));
assign main_rtio_core_inputs_blindtransfer7_i = main_rtio_core_inputs_overflow_io7;
assign main_rtio_core_inputs_selected7 = (main_rtio_core_cri_chan_sel[15:0] == 3'd7);
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_re = ((main_rtio_core_inputs_selected7 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow7));
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_din = {main_rtio_core_inputs_record8_fifo_in_data};
assign {main_rtio_core_inputs_record8_fifo_out_data} = main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout;
assign main_rtio_core_inputs_record8_fifo_in_data = main_spimaster0_iinterface0_data;
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_we = main_spimaster0_iinterface0_stb;
assign main_rtio_core_inputs_overflow_io8 = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_we & (~main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable));
assign main_rtio_core_inputs_blindtransfer8_i = main_rtio_core_inputs_overflow_io8;
assign main_rtio_core_inputs_selected8 = (main_rtio_core_cri_chan_sel[15:0] == 5'd16);
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_re = ((main_rtio_core_inputs_selected8 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow8));
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_din = {main_rtio_core_inputs_record9_fifo_in_data};
assign {main_rtio_core_inputs_record9_fifo_out_data} = main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout;
assign main_rtio_core_inputs_record9_fifo_in_data = main_spimaster1_iinterface1_data;
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_we = main_spimaster1_iinterface1_stb;
assign main_rtio_core_inputs_overflow_io9 = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_we & (~main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable));
assign main_rtio_core_inputs_blindtransfer9_i = main_rtio_core_inputs_overflow_io9;
assign main_rtio_core_inputs_selected9 = (main_rtio_core_cri_chan_sel[15:0] == 5'd22);
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_re = ((main_rtio_core_inputs_selected9 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow9));
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_din = {main_rtio_core_inputs_record10_fifo_in_data};
assign {main_rtio_core_inputs_record10_fifo_out_data} = main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout;
assign main_rtio_core_inputs_record10_fifo_in_data = main_spimaster2_iinterface2_data;
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_we = main_spimaster2_iinterface2_stb;
assign main_rtio_core_inputs_overflow_io10 = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_we & (~main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable));
assign main_rtio_core_inputs_blindtransfer10_i = main_rtio_core_inputs_overflow_io10;
assign main_rtio_core_inputs_selected10 = (main_rtio_core_cri_chan_sel[15:0] == 5'd28);
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_re = ((main_rtio_core_inputs_selected10 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow10));
assign main_rtio_core_inputs_i_status_raw = builder_comb_rhs_array_muxed9;
assign main_rtio_core_inputs_asyncfifo0_graycounter0_ce = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable & main_rtio_core_inputs_asyncfifo0_asyncfifo0_we);
assign main_rtio_core_inputs_asyncfifo0_graycounter1_ce = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & main_rtio_core_inputs_asyncfifo0_asyncfifo0_re);
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable = (((main_rtio_core_inputs_asyncfifo0_graycounter0_q[6] == main_rtio_core_inputs_asyncfifo0_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo0_graycounter0_q[5] == main_rtio_core_inputs_asyncfifo0_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo0_graycounter0_q[4:0] != main_rtio_core_inputs_asyncfifo0_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable = (main_rtio_core_inputs_asyncfifo0_graycounter1_q != main_rtio_core_inputs_asyncfifo0_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo0_wrport_adr = main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo0_wrport_dat_w = main_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
assign main_rtio_core_inputs_asyncfifo0_wrport_we = main_rtio_core_inputs_asyncfifo0_graycounter0_ce;
assign main_rtio_core_inputs_asyncfifo0_rdport_adr = main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout = main_rtio_core_inputs_asyncfifo0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_132;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo0_graycounter0_ce) begin
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= (main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_132 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_graycounter0_q_next = (main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary ^ main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_133;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo0_graycounter1_ce) begin
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= (main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_133 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_graycounter1_q_next = (main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary ^ main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer0_ps_i = (main_rtio_core_inputs_blindtransfer0_i & (~main_rtio_core_inputs_blindtransfer0_blind));
assign main_rtio_core_inputs_blindtransfer0_ps_ack_i = main_rtio_core_inputs_blindtransfer0_ps_o;
assign main_rtio_core_inputs_blindtransfer0_o = main_rtio_core_inputs_blindtransfer0_ps_o;
assign main_rtio_core_inputs_blindtransfer0_ps_o = (main_rtio_core_inputs_blindtransfer0_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer0_ps_ack_o = (main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo1_graycounter2_ce = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable & main_rtio_core_inputs_asyncfifo1_asyncfifo1_we);
assign main_rtio_core_inputs_asyncfifo1_graycounter3_ce = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & main_rtio_core_inputs_asyncfifo1_asyncfifo1_re);
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable = (((main_rtio_core_inputs_asyncfifo1_graycounter2_q[6] == main_rtio_core_inputs_asyncfifo1_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo1_graycounter2_q[5] == main_rtio_core_inputs_asyncfifo1_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo1_graycounter2_q[4:0] != main_rtio_core_inputs_asyncfifo1_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable = (main_rtio_core_inputs_asyncfifo1_graycounter3_q != main_rtio_core_inputs_asyncfifo1_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo1_wrport_adr = main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo1_wrport_dat_w = main_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
assign main_rtio_core_inputs_asyncfifo1_wrport_we = main_rtio_core_inputs_asyncfifo1_graycounter2_ce;
assign main_rtio_core_inputs_asyncfifo1_rdport_adr = main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout = main_rtio_core_inputs_asyncfifo1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_134;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo1_graycounter2_ce) begin
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= (main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_134 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo1_graycounter2_q_next = (main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary ^ main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_135;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo1_graycounter3_ce) begin
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= (main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_135 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo1_graycounter3_q_next = (main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary ^ main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer1_ps_i = (main_rtio_core_inputs_blindtransfer1_i & (~main_rtio_core_inputs_blindtransfer1_blind));
assign main_rtio_core_inputs_blindtransfer1_ps_ack_i = main_rtio_core_inputs_blindtransfer1_ps_o;
assign main_rtio_core_inputs_blindtransfer1_o = main_rtio_core_inputs_blindtransfer1_ps_o;
assign main_rtio_core_inputs_blindtransfer1_ps_o = (main_rtio_core_inputs_blindtransfer1_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer1_ps_ack_o = (main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo2_graycounter4_ce = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable & main_rtio_core_inputs_asyncfifo2_asyncfifo2_we);
assign main_rtio_core_inputs_asyncfifo2_graycounter5_ce = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & main_rtio_core_inputs_asyncfifo2_asyncfifo2_re);
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable = (((main_rtio_core_inputs_asyncfifo2_graycounter4_q[6] == main_rtio_core_inputs_asyncfifo2_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo2_graycounter4_q[5] == main_rtio_core_inputs_asyncfifo2_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo2_graycounter4_q[4:0] != main_rtio_core_inputs_asyncfifo2_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable = (main_rtio_core_inputs_asyncfifo2_graycounter5_q != main_rtio_core_inputs_asyncfifo2_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo2_wrport_adr = main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo2_wrport_dat_w = main_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
assign main_rtio_core_inputs_asyncfifo2_wrport_we = main_rtio_core_inputs_asyncfifo2_graycounter4_ce;
assign main_rtio_core_inputs_asyncfifo2_rdport_adr = main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout = main_rtio_core_inputs_asyncfifo2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_136;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo2_graycounter4_ce) begin
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= (main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_136 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo2_graycounter4_q_next = (main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary ^ main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_137;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo2_graycounter5_ce) begin
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= (main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_137 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo2_graycounter5_q_next = (main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary ^ main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer2_ps_i = (main_rtio_core_inputs_blindtransfer2_i & (~main_rtio_core_inputs_blindtransfer2_blind));
assign main_rtio_core_inputs_blindtransfer2_ps_ack_i = main_rtio_core_inputs_blindtransfer2_ps_o;
assign main_rtio_core_inputs_blindtransfer2_o = main_rtio_core_inputs_blindtransfer2_ps_o;
assign main_rtio_core_inputs_blindtransfer2_ps_o = (main_rtio_core_inputs_blindtransfer2_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer2_ps_ack_o = (main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo3_graycounter6_ce = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable & main_rtio_core_inputs_asyncfifo3_asyncfifo3_we);
assign main_rtio_core_inputs_asyncfifo3_graycounter7_ce = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & main_rtio_core_inputs_asyncfifo3_asyncfifo3_re);
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable = (((main_rtio_core_inputs_asyncfifo3_graycounter6_q[6] == main_rtio_core_inputs_asyncfifo3_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo3_graycounter6_q[5] == main_rtio_core_inputs_asyncfifo3_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo3_graycounter6_q[4:0] != main_rtio_core_inputs_asyncfifo3_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable = (main_rtio_core_inputs_asyncfifo3_graycounter7_q != main_rtio_core_inputs_asyncfifo3_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo3_wrport_adr = main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo3_wrport_dat_w = main_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
assign main_rtio_core_inputs_asyncfifo3_wrport_we = main_rtio_core_inputs_asyncfifo3_graycounter6_ce;
assign main_rtio_core_inputs_asyncfifo3_rdport_adr = main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout = main_rtio_core_inputs_asyncfifo3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_138;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo3_graycounter6_ce) begin
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= (main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_138 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo3_graycounter6_q_next = (main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary ^ main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_139;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo3_graycounter7_ce) begin
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= (main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_139 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo3_graycounter7_q_next = (main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary ^ main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer3_ps_i = (main_rtio_core_inputs_blindtransfer3_i & (~main_rtio_core_inputs_blindtransfer3_blind));
assign main_rtio_core_inputs_blindtransfer3_ps_ack_i = main_rtio_core_inputs_blindtransfer3_ps_o;
assign main_rtio_core_inputs_blindtransfer3_o = main_rtio_core_inputs_blindtransfer3_ps_o;
assign main_rtio_core_inputs_blindtransfer3_ps_o = (main_rtio_core_inputs_blindtransfer3_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer3_ps_ack_o = (main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo4_graycounter8_ce = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable & main_rtio_core_inputs_asyncfifo4_asyncfifo4_we);
assign main_rtio_core_inputs_asyncfifo4_graycounter9_ce = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & main_rtio_core_inputs_asyncfifo4_asyncfifo4_re);
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable = (((main_rtio_core_inputs_asyncfifo4_graycounter8_q[6] == main_rtio_core_inputs_asyncfifo4_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo4_graycounter8_q[5] == main_rtio_core_inputs_asyncfifo4_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo4_graycounter8_q[4:0] != main_rtio_core_inputs_asyncfifo4_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable = (main_rtio_core_inputs_asyncfifo4_graycounter9_q != main_rtio_core_inputs_asyncfifo4_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo4_wrport_adr = main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo4_wrport_dat_w = main_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
assign main_rtio_core_inputs_asyncfifo4_wrport_we = main_rtio_core_inputs_asyncfifo4_graycounter8_ce;
assign main_rtio_core_inputs_asyncfifo4_rdport_adr = main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout = main_rtio_core_inputs_asyncfifo4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_140;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo4_graycounter8_ce) begin
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= (main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_140 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo4_graycounter8_q_next = (main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary ^ main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_141;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo4_graycounter9_ce) begin
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= (main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_141 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo4_graycounter9_q_next = (main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary ^ main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer4_ps_i = (main_rtio_core_inputs_blindtransfer4_i & (~main_rtio_core_inputs_blindtransfer4_blind));
assign main_rtio_core_inputs_blindtransfer4_ps_ack_i = main_rtio_core_inputs_blindtransfer4_ps_o;
assign main_rtio_core_inputs_blindtransfer4_o = main_rtio_core_inputs_blindtransfer4_ps_o;
assign main_rtio_core_inputs_blindtransfer4_ps_o = (main_rtio_core_inputs_blindtransfer4_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer4_ps_ack_o = (main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo5_graycounter10_ce = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable & main_rtio_core_inputs_asyncfifo5_asyncfifo5_we);
assign main_rtio_core_inputs_asyncfifo5_graycounter11_ce = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & main_rtio_core_inputs_asyncfifo5_asyncfifo5_re);
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable = (((main_rtio_core_inputs_asyncfifo5_graycounter10_q[6] == main_rtio_core_inputs_asyncfifo5_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo5_graycounter10_q[5] == main_rtio_core_inputs_asyncfifo5_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo5_graycounter10_q[4:0] != main_rtio_core_inputs_asyncfifo5_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable = (main_rtio_core_inputs_asyncfifo5_graycounter11_q != main_rtio_core_inputs_asyncfifo5_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo5_wrport_adr = main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo5_wrport_dat_w = main_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
assign main_rtio_core_inputs_asyncfifo5_wrport_we = main_rtio_core_inputs_asyncfifo5_graycounter10_ce;
assign main_rtio_core_inputs_asyncfifo5_rdport_adr = main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout = main_rtio_core_inputs_asyncfifo5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_142;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo5_graycounter10_ce) begin
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= (main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_142 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo5_graycounter10_q_next = (main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary ^ main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_143;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo5_graycounter11_ce) begin
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= (main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_143 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo5_graycounter11_q_next = (main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary ^ main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer5_ps_i = (main_rtio_core_inputs_blindtransfer5_i & (~main_rtio_core_inputs_blindtransfer5_blind));
assign main_rtio_core_inputs_blindtransfer5_ps_ack_i = main_rtio_core_inputs_blindtransfer5_ps_o;
assign main_rtio_core_inputs_blindtransfer5_o = main_rtio_core_inputs_blindtransfer5_ps_o;
assign main_rtio_core_inputs_blindtransfer5_ps_o = (main_rtio_core_inputs_blindtransfer5_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer5_ps_ack_o = (main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo6_graycounter12_ce = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable & main_rtio_core_inputs_asyncfifo6_asyncfifo6_we);
assign main_rtio_core_inputs_asyncfifo6_graycounter13_ce = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & main_rtio_core_inputs_asyncfifo6_asyncfifo6_re);
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable = (((main_rtio_core_inputs_asyncfifo6_graycounter12_q[6] == main_rtio_core_inputs_asyncfifo6_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo6_graycounter12_q[5] == main_rtio_core_inputs_asyncfifo6_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo6_graycounter12_q[4:0] != main_rtio_core_inputs_asyncfifo6_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable = (main_rtio_core_inputs_asyncfifo6_graycounter13_q != main_rtio_core_inputs_asyncfifo6_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo6_wrport_adr = main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo6_wrport_dat_w = main_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
assign main_rtio_core_inputs_asyncfifo6_wrport_we = main_rtio_core_inputs_asyncfifo6_graycounter12_ce;
assign main_rtio_core_inputs_asyncfifo6_rdport_adr = main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout = main_rtio_core_inputs_asyncfifo6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_144;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo6_graycounter12_ce) begin
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= (main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_144 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo6_graycounter12_q_next = (main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary ^ main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_145;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo6_graycounter13_ce) begin
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= (main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_145 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo6_graycounter13_q_next = (main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary ^ main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer6_ps_i = (main_rtio_core_inputs_blindtransfer6_i & (~main_rtio_core_inputs_blindtransfer6_blind));
assign main_rtio_core_inputs_blindtransfer6_ps_ack_i = main_rtio_core_inputs_blindtransfer6_ps_o;
assign main_rtio_core_inputs_blindtransfer6_o = main_rtio_core_inputs_blindtransfer6_ps_o;
assign main_rtio_core_inputs_blindtransfer6_ps_o = (main_rtio_core_inputs_blindtransfer6_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer6_ps_ack_o = (main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo7_graycounter14_ce = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable & main_rtio_core_inputs_asyncfifo7_asyncfifo7_we);
assign main_rtio_core_inputs_asyncfifo7_graycounter15_ce = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable & main_rtio_core_inputs_asyncfifo7_asyncfifo7_re);
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable = (((main_rtio_core_inputs_asyncfifo7_graycounter14_q[6] == main_rtio_core_inputs_asyncfifo7_consume_wdomain[6]) | (main_rtio_core_inputs_asyncfifo7_graycounter14_q[5] == main_rtio_core_inputs_asyncfifo7_consume_wdomain[5])) | (main_rtio_core_inputs_asyncfifo7_graycounter14_q[4:0] != main_rtio_core_inputs_asyncfifo7_consume_wdomain[4:0]));
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable = (main_rtio_core_inputs_asyncfifo7_graycounter15_q != main_rtio_core_inputs_asyncfifo7_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo7_wrport_adr = main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary[5:0];
assign main_rtio_core_inputs_asyncfifo7_wrport_dat_w = main_rtio_core_inputs_asyncfifo7_asyncfifo7_din;
assign main_rtio_core_inputs_asyncfifo7_wrport_we = main_rtio_core_inputs_asyncfifo7_graycounter14_ce;
assign main_rtio_core_inputs_asyncfifo7_rdport_adr = main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary[5:0];
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout = main_rtio_core_inputs_asyncfifo7_rdport_dat_r;

// synthesis translate_off
reg dummy_d_146;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo7_graycounter14_ce) begin
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= (main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary;
	end
// synthesis translate_off
	dummy_d_146 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo7_graycounter14_q_next = (main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary ^ main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_147;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= 7'd0;
	if (main_rtio_core_inputs_asyncfifo7_graycounter15_ce) begin
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= (main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary;
	end
// synthesis translate_off
	dummy_d_147 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo7_graycounter15_q_next = (main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary ^ main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary[6:1]);
assign main_rtio_core_inputs_blindtransfer7_ps_i = (main_rtio_core_inputs_blindtransfer7_i & (~main_rtio_core_inputs_blindtransfer7_blind));
assign main_rtio_core_inputs_blindtransfer7_ps_ack_i = main_rtio_core_inputs_blindtransfer7_ps_o;
assign main_rtio_core_inputs_blindtransfer7_o = main_rtio_core_inputs_blindtransfer7_ps_o;
assign main_rtio_core_inputs_blindtransfer7_ps_o = (main_rtio_core_inputs_blindtransfer7_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer7_ps_ack_o = (main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo8_graycounter16_ce = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable & main_rtio_core_inputs_asyncfifo8_asyncfifo8_we);
assign main_rtio_core_inputs_asyncfifo8_graycounter17_ce = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable & main_rtio_core_inputs_asyncfifo8_asyncfifo8_re);
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable = (((main_rtio_core_inputs_asyncfifo8_graycounter16_q[2] == main_rtio_core_inputs_asyncfifo8_consume_wdomain[2]) | (main_rtio_core_inputs_asyncfifo8_graycounter16_q[1] == main_rtio_core_inputs_asyncfifo8_consume_wdomain[1])) | (main_rtio_core_inputs_asyncfifo8_graycounter16_q[0] != main_rtio_core_inputs_asyncfifo8_consume_wdomain[0]));
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable = (main_rtio_core_inputs_asyncfifo8_graycounter17_q != main_rtio_core_inputs_asyncfifo8_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo8_wrport_adr = main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary[1:0];
assign main_rtio_core_inputs_asyncfifo8_wrport_dat_w = main_rtio_core_inputs_asyncfifo8_asyncfifo8_din;
assign main_rtio_core_inputs_asyncfifo8_wrport_we = main_rtio_core_inputs_asyncfifo8_graycounter16_ce;
assign main_rtio_core_inputs_asyncfifo8_rdport_adr = main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary[1:0];
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout = main_rtio_core_inputs_asyncfifo8_rdport_dat_r;

// synthesis translate_off
reg dummy_d_148;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo8_graycounter16_ce) begin
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= (main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary;
	end
// synthesis translate_off
	dummy_d_148 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo8_graycounter16_q_next = (main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary ^ main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_149;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo8_graycounter17_ce) begin
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= (main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary;
	end
// synthesis translate_off
	dummy_d_149 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo8_graycounter17_q_next = (main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary ^ main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary[2:1]);
assign main_rtio_core_inputs_blindtransfer8_ps_i = (main_rtio_core_inputs_blindtransfer8_i & (~main_rtio_core_inputs_blindtransfer8_blind));
assign main_rtio_core_inputs_blindtransfer8_ps_ack_i = main_rtio_core_inputs_blindtransfer8_ps_o;
assign main_rtio_core_inputs_blindtransfer8_o = main_rtio_core_inputs_blindtransfer8_ps_o;
assign main_rtio_core_inputs_blindtransfer8_ps_o = (main_rtio_core_inputs_blindtransfer8_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer8_ps_ack_o = (main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo9_graycounter18_ce = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable & main_rtio_core_inputs_asyncfifo9_asyncfifo9_we);
assign main_rtio_core_inputs_asyncfifo9_graycounter19_ce = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable & main_rtio_core_inputs_asyncfifo9_asyncfifo9_re);
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable = (((main_rtio_core_inputs_asyncfifo9_graycounter18_q[2] == main_rtio_core_inputs_asyncfifo9_consume_wdomain[2]) | (main_rtio_core_inputs_asyncfifo9_graycounter18_q[1] == main_rtio_core_inputs_asyncfifo9_consume_wdomain[1])) | (main_rtio_core_inputs_asyncfifo9_graycounter18_q[0] != main_rtio_core_inputs_asyncfifo9_consume_wdomain[0]));
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable = (main_rtio_core_inputs_asyncfifo9_graycounter19_q != main_rtio_core_inputs_asyncfifo9_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo9_wrport_adr = main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary[1:0];
assign main_rtio_core_inputs_asyncfifo9_wrport_dat_w = main_rtio_core_inputs_asyncfifo9_asyncfifo9_din;
assign main_rtio_core_inputs_asyncfifo9_wrport_we = main_rtio_core_inputs_asyncfifo9_graycounter18_ce;
assign main_rtio_core_inputs_asyncfifo9_rdport_adr = main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary[1:0];
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout = main_rtio_core_inputs_asyncfifo9_rdport_dat_r;

// synthesis translate_off
reg dummy_d_150;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo9_graycounter18_ce) begin
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= (main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary;
	end
// synthesis translate_off
	dummy_d_150 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo9_graycounter18_q_next = (main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary ^ main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_151;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo9_graycounter19_ce) begin
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= (main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary;
	end
// synthesis translate_off
	dummy_d_151 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo9_graycounter19_q_next = (main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary ^ main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary[2:1]);
assign main_rtio_core_inputs_blindtransfer9_ps_i = (main_rtio_core_inputs_blindtransfer9_i & (~main_rtio_core_inputs_blindtransfer9_blind));
assign main_rtio_core_inputs_blindtransfer9_ps_ack_i = main_rtio_core_inputs_blindtransfer9_ps_o;
assign main_rtio_core_inputs_blindtransfer9_o = main_rtio_core_inputs_blindtransfer9_ps_o;
assign main_rtio_core_inputs_blindtransfer9_ps_o = (main_rtio_core_inputs_blindtransfer9_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer9_ps_ack_o = (main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo10_graycounter20_ce = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable & main_rtio_core_inputs_asyncfifo10_asyncfifo10_we);
assign main_rtio_core_inputs_asyncfifo10_graycounter21_ce = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable & main_rtio_core_inputs_asyncfifo10_asyncfifo10_re);
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable = (((main_rtio_core_inputs_asyncfifo10_graycounter20_q[2] == main_rtio_core_inputs_asyncfifo10_consume_wdomain[2]) | (main_rtio_core_inputs_asyncfifo10_graycounter20_q[1] == main_rtio_core_inputs_asyncfifo10_consume_wdomain[1])) | (main_rtio_core_inputs_asyncfifo10_graycounter20_q[0] != main_rtio_core_inputs_asyncfifo10_consume_wdomain[0]));
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable = (main_rtio_core_inputs_asyncfifo10_graycounter21_q != main_rtio_core_inputs_asyncfifo10_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo10_wrport_adr = main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary[1:0];
assign main_rtio_core_inputs_asyncfifo10_wrport_dat_w = main_rtio_core_inputs_asyncfifo10_asyncfifo10_din;
assign main_rtio_core_inputs_asyncfifo10_wrport_we = main_rtio_core_inputs_asyncfifo10_graycounter20_ce;
assign main_rtio_core_inputs_asyncfifo10_rdport_adr = main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary[1:0];
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout = main_rtio_core_inputs_asyncfifo10_rdport_dat_r;

// synthesis translate_off
reg dummy_d_152;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo10_graycounter20_ce) begin
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= (main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary;
	end
// synthesis translate_off
	dummy_d_152 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo10_graycounter20_q_next = (main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary ^ main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_153;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo10_graycounter21_ce) begin
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= (main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary;
	end
// synthesis translate_off
	dummy_d_153 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo10_graycounter21_q_next = (main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary ^ main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary[2:1]);
assign main_rtio_core_inputs_blindtransfer10_ps_i = (main_rtio_core_inputs_blindtransfer10_i & (~main_rtio_core_inputs_blindtransfer10_blind));
assign main_rtio_core_inputs_blindtransfer10_ps_ack_i = main_rtio_core_inputs_blindtransfer10_ps_o;
assign main_rtio_core_inputs_blindtransfer10_o = main_rtio_core_inputs_blindtransfer10_ps_o;
assign main_rtio_core_inputs_blindtransfer10_ps_o = (main_rtio_core_inputs_blindtransfer10_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer10_ps_ack_o = (main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r);
assign main_rtio_core_o_collision_sync_ps_i = (main_rtio_core_o_collision_sync_i & (~main_rtio_core_o_collision_sync_blind));
assign main_rtio_core_o_collision_sync_ps_ack_i = main_rtio_core_o_collision_sync_ps_o;
assign main_rtio_core_o_collision_sync_o = main_rtio_core_o_collision_sync_ps_o;
assign main_rtio_core_o_collision_sync_ps_o = (main_rtio_core_o_collision_sync_ps_toggle_o ^ main_rtio_core_o_collision_sync_ps_toggle_o_r);
assign main_rtio_core_o_collision_sync_ps_ack_o = (main_rtio_core_o_collision_sync_ps_ack_toggle_o ^ main_rtio_core_o_collision_sync_ps_ack_toggle_o_r);
assign main_rtio_core_o_busy_sync_ps_i = (main_rtio_core_o_busy_sync_i & (~main_rtio_core_o_busy_sync_blind));
assign main_rtio_core_o_busy_sync_ps_ack_i = main_rtio_core_o_busy_sync_ps_o;
assign main_rtio_core_o_busy_sync_o = main_rtio_core_o_busy_sync_ps_o;
assign main_rtio_core_o_busy_sync_ps_o = (main_rtio_core_o_busy_sync_ps_toggle_o ^ main_rtio_core_o_busy_sync_ps_toggle_o_r);
assign main_rtio_core_o_busy_sync_ps_ack_o = (main_rtio_core_o_busy_sync_ps_ack_toggle_o ^ main_rtio_core_o_busy_sync_ps_ack_toggle_o_r);
assign main_rtio_now_hi_w = main_rtio_now[63:32];
assign main_rtio_now_lo_w = main_rtio_now[31:0];

// synthesis translate_off
reg dummy_d_154;
// synthesis translate_on
always @(*) begin
	main_rtio_cri_cmd <= 2'd0;
	main_rtio_cri_cmd <= 1'd0;
	if (main_rtio_o_data_re) begin
		main_rtio_cri_cmd <= 1'd1;
	end
	if (main_rtio_i_timeout_re) begin
		main_rtio_cri_cmd <= 2'd2;
	end
// synthesis translate_off
	dummy_d_154 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_cri_chan_sel = main_rtio_target_storage[31:8];
assign main_rtio_cri_o_timestamp = main_rtio_now;
assign main_rtio_cri_o_data = main_rtio_o_data_storage;
assign main_rtio_cri_o_address = main_rtio_target_storage[7:0];
assign main_rtio_o_status_status = main_rtio_cri_o_status;
assign main_rtio_cri_i_timeout = main_rtio_i_timeout_storage;
assign main_rtio_i_data_status = main_rtio_cri_i_data;
assign main_rtio_i_timestamp_status = main_rtio_cri_i_timestamp;
assign main_rtio_i_status_status = main_rtio_cri_i_status;
assign main_rtio_o_data_dat_w = 1'd0;
assign main_rtio_o_data_we = main_rtio_target_re;
assign main_dma_rawslicer_sink_stb = main_dma_dma_source_stb;
assign main_dma_dma_source_ack = main_dma_rawslicer_sink_ack;
assign main_dma_rawslicer_sink_eop = main_dma_dma_source_eop;
assign main_dma_rawslicer_sink_payload_data = main_dma_dma_source_payload_data;
assign main_dma_time_offset_sink_stb = main_dma_record_converter_source_stb;
assign main_dma_record_converter_source_ack = main_dma_time_offset_sink_ack;
assign main_dma_time_offset_sink_eop = main_dma_record_converter_source_eop;
assign main_dma_time_offset_sink_payload_length = main_dma_record_converter_source_payload_length;
assign main_dma_time_offset_sink_payload_channel = main_dma_record_converter_source_payload_channel;
assign main_dma_time_offset_sink_payload_timestamp = main_dma_record_converter_source_payload_timestamp;
assign main_dma_time_offset_sink_payload_address = main_dma_record_converter_source_payload_address;
assign main_dma_time_offset_sink_payload_data = main_dma_record_converter_source_payload_data;
assign main_dma_cri_master_sink_stb = main_dma_time_offset_source_stb;
assign main_dma_time_offset_source_ack = main_dma_cri_master_sink_ack;
assign main_dma_cri_master_sink_eop = main_dma_time_offset_source_eop;
assign main_dma_cri_master_sink_payload_length = main_dma_time_offset_source_payload_length;
assign main_dma_cri_master_sink_payload_channel = main_dma_time_offset_source_payload_channel;
assign main_dma_cri_master_sink_payload_timestamp = main_dma_time_offset_source_payload_timestamp;
assign main_dma_cri_master_sink_payload_address = main_dma_time_offset_source_payload_address;
assign main_dma_cri_master_sink_payload_data = main_dma_time_offset_source_payload_data;
assign main_dma_dma_bus_stb = (main_dma_dma_sink_stb & ((~main_dma_dma_data_reg_loaded) | main_dma_dma_source_ack));
assign main_genericstandalone_interface0_bus_cyc = main_dma_dma_bus_stb;
assign main_genericstandalone_interface0_bus_stb = main_dma_dma_bus_stb;
assign main_genericstandalone_interface0_bus_adr = main_dma_dma_sink_payload_address;
assign main_dma_dma_sink_ack = main_genericstandalone_interface0_bus_ack;
assign main_dma_dma_source_stb = main_dma_dma_data_reg_loaded;
assign main_dma_rawslicer_source = main_dma_rawslicer_buf[615:0];

// synthesis translate_off
reg dummy_d_155;
// synthesis translate_on
always @(*) begin
	main_dma_rawslicer_sink_ack <= 1'd0;
	main_dma_rawslicer_source_stb <= 1'd0;
	main_dma_rawslicer_flush_done <= 1'd0;
	main_dma_rawslicer_next_level <= 7'd0;
	main_dma_rawslicer_load_buf <= 1'd0;
	main_dma_rawslicer_shift_buf <= 1'd0;
	builder_clockdomainsrenamer_resetinserter_next_state <= 2'd0;
	main_dma_rawslicer_next_level <= main_dma_rawslicer_level;
	builder_clockdomainsrenamer_resetinserter_next_state <= builder_clockdomainsrenamer_resetinserter_state;
	case (builder_clockdomainsrenamer_resetinserter_state)
		1'd1: begin
			main_dma_rawslicer_source_stb <= 1'd1;
			main_dma_rawslicer_shift_buf <= 1'd1;
			main_dma_rawslicer_next_level <= (main_dma_rawslicer_level - main_dma_rawslicer_source_consume);
			if ((main_dma_rawslicer_next_level < 7'd77)) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
			if (main_dma_rawslicer_flush) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_dma_rawslicer_next_level <= 1'd0;
			main_dma_rawslicer_sink_ack <= 1'd1;
			if ((main_dma_rawslicer_sink_stb & main_dma_rawslicer_sink_eop)) begin
				main_dma_rawslicer_flush_done <= 1'd1;
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_dma_rawslicer_sink_ack <= 1'd1;
			main_dma_rawslicer_load_buf <= 1'd1;
			if (main_dma_rawslicer_sink_stb) begin
				main_dma_rawslicer_next_level <= (main_dma_rawslicer_level + 5'd16);
			end
			if ((main_dma_rawslicer_next_level >= 7'd77)) begin
				builder_clockdomainsrenamer_resetinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_155 <= dummy_s;
// synthesis translate_on
end
assign {main_dma_record_converter_record_raw_data, main_dma_record_converter_record_raw_address, main_dma_record_converter_record_raw_timestamp, main_dma_record_converter_record_raw_channel, main_dma_record_converter_record_raw_length} = main_dma_rawslicer_source;
assign main_dma_record_converter_source_payload_channel = main_dma_record_converter_record_raw_channel;
assign main_dma_record_converter_source_payload_timestamp = main_dma_record_converter_record_raw_timestamp;
assign main_dma_record_converter_source_payload_address = main_dma_record_converter_record_raw_address;

// synthesis translate_off
reg dummy_d_156;
// synthesis translate_on
always @(*) begin
	main_dma_record_converter_source_payload_data <= 512'd0;
	case (main_dma_record_converter_record_raw_length)
		4'd14: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[7:0];
		end
		4'd15: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[15:0];
		end
		5'd16: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[23:0];
		end
		5'd17: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[31:0];
		end
		5'd18: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[39:0];
		end
		5'd19: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[47:0];
		end
		5'd20: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[55:0];
		end
		5'd21: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[63:0];
		end
		5'd22: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[71:0];
		end
		5'd23: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[79:0];
		end
		5'd24: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[87:0];
		end
		5'd25: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[95:0];
		end
		5'd26: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[103:0];
		end
		5'd27: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[111:0];
		end
		5'd28: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[119:0];
		end
		5'd29: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[127:0];
		end
		5'd30: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[135:0];
		end
		5'd31: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[143:0];
		end
		6'd32: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[151:0];
		end
		6'd33: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[159:0];
		end
		6'd34: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[167:0];
		end
		6'd35: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[175:0];
		end
		6'd36: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[183:0];
		end
		6'd37: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[191:0];
		end
		6'd38: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[199:0];
		end
		6'd39: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[207:0];
		end
		6'd40: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[215:0];
		end
		6'd41: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[223:0];
		end
		6'd42: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[231:0];
		end
		6'd43: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[239:0];
		end
		6'd44: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[247:0];
		end
		6'd45: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[255:0];
		end
		6'd46: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[263:0];
		end
		6'd47: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[271:0];
		end
		6'd48: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[279:0];
		end
		6'd49: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[287:0];
		end
		6'd50: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[295:0];
		end
		6'd51: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[303:0];
		end
		6'd52: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[311:0];
		end
		6'd53: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[319:0];
		end
		6'd54: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[327:0];
		end
		6'd55: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[335:0];
		end
		6'd56: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[343:0];
		end
		6'd57: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[351:0];
		end
		6'd58: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[359:0];
		end
		6'd59: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[367:0];
		end
		6'd60: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[375:0];
		end
		6'd61: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[383:0];
		end
		6'd62: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[391:0];
		end
		6'd63: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[399:0];
		end
		7'd64: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[407:0];
		end
		7'd65: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[415:0];
		end
		7'd66: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[423:0];
		end
		7'd67: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[431:0];
		end
		7'd68: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[439:0];
		end
		7'd69: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[447:0];
		end
		7'd70: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[455:0];
		end
		7'd71: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[463:0];
		end
		7'd72: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[471:0];
		end
		7'd73: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[479:0];
		end
		7'd74: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[487:0];
		end
		7'd75: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[495:0];
		end
		7'd76: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[503:0];
		end
		7'd77: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[511:0];
		end
	endcase
// synthesis translate_off
	dummy_d_156 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_157;
// synthesis translate_on
always @(*) begin
	main_dma_rawslicer_source_consume <= 7'd0;
	main_dma_rawslicer_flush <= 1'd0;
	main_dma_record_converter_source_stb <= 1'd0;
	main_dma_record_converter_source_eop <= 1'd0;
	main_dma_record_converter_end_marker_found <= 1'd0;
	builder_clockdomainsrenamer_recordconverter_next_state <= 2'd0;
	builder_clockdomainsrenamer_recordconverter_next_state <= builder_clockdomainsrenamer_recordconverter_state;
	case (builder_clockdomainsrenamer_recordconverter_state)
		1'd1: begin
			main_dma_record_converter_end_marker_found <= 1'd1;
			if (main_dma_record_converter_flush) begin
				main_dma_rawslicer_flush <= 1'd1;
				builder_clockdomainsrenamer_recordconverter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (main_dma_rawslicer_flush_done) begin
				builder_clockdomainsrenamer_recordconverter_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_dma_record_converter_source_eop <= 1'd1;
			main_dma_record_converter_source_stb <= 1'd1;
			if (main_dma_record_converter_source_ack) begin
				builder_clockdomainsrenamer_recordconverter_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_dma_rawslicer_source_stb) begin
				if ((main_dma_record_converter_record_raw_length == 1'd0)) begin
					builder_clockdomainsrenamer_recordconverter_next_state <= 1'd1;
				end else begin
					main_dma_record_converter_source_stb <= 1'd1;
				end
			end
			if (main_dma_record_converter_source_ack) begin
				main_dma_rawslicer_source_consume <= main_dma_record_converter_record_raw_length;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_157 <= dummy_s;
// synthesis translate_on
end
assign main_dma_time_offset_sink_ack = (~main_dma_time_offset_source_stb);
assign main_dma_cri_master_cri_chan_sel = main_dma_cri_master_sink_payload_channel;
assign main_dma_cri_master_cri_o_timestamp = main_dma_cri_master_sink_payload_timestamp;
assign main_dma_cri_master_cri_o_address = main_dma_cri_master_sink_payload_address;
assign main_dma_cri_master_cri_o_data = main_dma_cri_master_sink_payload_data;

// synthesis translate_off
reg dummy_d_158;
// synthesis translate_on
always @(*) begin
	main_dma_cri_master_sink_ack <= 1'd0;
	main_dma_cri_master_cri_cmd <= 2'd0;
	main_dma_cri_master_busy <= 1'd0;
	main_dma_cri_master_underflow_trigger <= 1'd0;
	main_dma_cri_master_link_error_trigger <= 1'd0;
	builder_clockdomainsrenamer_crimaster_next_state <= 3'd0;
	builder_clockdomainsrenamer_crimaster_next_state <= builder_clockdomainsrenamer_crimaster_state;
	case (builder_clockdomainsrenamer_crimaster_state)
		1'd1: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_cri_cmd <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 2'd2;
		end
		2'd2: begin
			main_dma_cri_master_busy <= 1'd1;
			if ((main_dma_cri_master_cri_o_status == 1'd0)) begin
				main_dma_cri_master_sink_ack <= 1'd1;
				builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
			end
			if (main_dma_cri_master_cri_o_status[1]) begin
				builder_clockdomainsrenamer_crimaster_next_state <= 2'd3;
			end
			if (main_dma_cri_master_cri_o_status[2]) begin
				builder_clockdomainsrenamer_crimaster_next_state <= 3'd4;
			end
		end
		2'd3: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_underflow_trigger <= 1'd1;
			main_dma_cri_master_sink_ack <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		3'd4: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_link_error_trigger <= 1'd1;
			main_dma_cri_master_sink_ack <= 1'd1;
			builder_clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		default: begin
			if ((main_dma_cri_master_error_w == 1'd0)) begin
				if (main_dma_cri_master_sink_stb) begin
					if (main_dma_cri_master_sink_eop) begin
						main_dma_cri_master_sink_ack <= 1'd1;
					end else begin
						builder_clockdomainsrenamer_crimaster_next_state <= 1'd1;
					end
				end
			end else begin
				main_dma_cri_master_sink_ack <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_158 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_159;
// synthesis translate_on
always @(*) begin
	main_dma_enable_enable_w <= 1'd0;
	main_dma_flow_enable <= 1'd0;
	main_dma_record_converter_flush <= 1'd0;
	builder_clockdomainsrenamer_fsm_next_state <= 3'd0;
	builder_clockdomainsrenamer_fsm_next_state <= builder_clockdomainsrenamer_fsm_state;
	case (builder_clockdomainsrenamer_fsm_state)
		1'd1: begin
			main_dma_enable_enable_w <= 1'd1;
			main_dma_flow_enable <= 1'd1;
			if (main_dma_record_converter_end_marker_found) begin
				builder_clockdomainsrenamer_fsm_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_dma_enable_enable_w <= 1'd1;
			main_dma_record_converter_flush <= 1'd1;
			builder_clockdomainsrenamer_fsm_next_state <= 2'd3;
		end
		2'd3: begin
			main_dma_enable_enable_w <= 1'd1;
			if (((main_dma_cri_master_sink_stb & main_dma_cri_master_sink_ack) & main_dma_cri_master_sink_eop)) begin
				builder_clockdomainsrenamer_fsm_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_dma_enable_enable_w <= 1'd1;
			if ((~main_dma_cri_master_busy)) begin
				builder_clockdomainsrenamer_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_dma_enable_enable_re) begin
				builder_clockdomainsrenamer_fsm_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_159 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_csrbank0_target0_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_target0_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 1'd0));
assign main_rtio_now_hi_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_rtio_now_hi_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 1'd1));
assign main_rtio_now_lo_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_rtio_now_lo_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 2'd2));
assign main_genericstandalone_csrbank0_o_data15_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data15_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 2'd3));
assign main_genericstandalone_csrbank0_o_data14_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data14_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 3'd4));
assign main_genericstandalone_csrbank0_o_data13_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data13_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 3'd5));
assign main_genericstandalone_csrbank0_o_data12_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data12_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 3'd6));
assign main_genericstandalone_csrbank0_o_data11_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data11_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 3'd7));
assign main_genericstandalone_csrbank0_o_data10_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data10_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd8));
assign main_genericstandalone_csrbank0_o_data9_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data9_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd9));
assign main_genericstandalone_csrbank0_o_data8_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data8_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd10));
assign main_genericstandalone_csrbank0_o_data7_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data7_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd11));
assign main_genericstandalone_csrbank0_o_data6_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data6_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd12));
assign main_genericstandalone_csrbank0_o_data5_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data5_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd13));
assign main_genericstandalone_csrbank0_o_data4_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data4_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd14));
assign main_genericstandalone_csrbank0_o_data3_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data3_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 4'd15));
assign main_genericstandalone_csrbank0_o_data2_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data2_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd16));
assign main_genericstandalone_csrbank0_o_data1_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data1_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd17));
assign main_genericstandalone_csrbank0_o_data0_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_o_data0_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd18));
assign main_genericstandalone_csrbank0_o_status_r = main_genericstandalone_csrbank0_bus_dat_w[2:0];
assign main_genericstandalone_csrbank0_o_status_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd19));
assign main_genericstandalone_csrbank0_i_timeout1_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_i_timeout1_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd20));
assign main_genericstandalone_csrbank0_i_timeout0_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_i_timeout0_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd21));
assign main_genericstandalone_csrbank0_i_data_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_i_data_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd22));
assign main_genericstandalone_csrbank0_i_timestamp1_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_i_timestamp1_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd23));
assign main_genericstandalone_csrbank0_i_timestamp0_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_i_timestamp0_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd24));
assign main_genericstandalone_csrbank0_i_status_r = main_genericstandalone_csrbank0_bus_dat_w[3:0];
assign main_genericstandalone_csrbank0_i_status_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd25));
assign main_rtio_i_overflow_reset_r = main_genericstandalone_csrbank0_bus_dat_w[0];
assign main_rtio_i_overflow_reset_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd26));
assign main_genericstandalone_csrbank0_counter1_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_counter1_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd27));
assign main_genericstandalone_csrbank0_counter0_r = main_genericstandalone_csrbank0_bus_dat_w[31:0];
assign main_genericstandalone_csrbank0_counter0_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd28));
assign main_rtio_counter_update_r = main_genericstandalone_csrbank0_bus_dat_w[0];
assign main_rtio_counter_update_re = ((((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb) & (~main_genericstandalone_csrbank0_bus_ack)) & main_genericstandalone_csrbank0_bus_we) & (main_genericstandalone_csrbank0_bus_adr[4:0] == 5'd29));
assign main_rtio_target_storage = main_rtio_target_storage_full[31:0];
assign main_genericstandalone_csrbank0_target0_w = main_rtio_target_storage_full[31:0];
assign main_rtio_o_data_storage = main_rtio_o_data_storage_full[511:0];
assign main_genericstandalone_csrbank0_o_data15_w = main_rtio_o_data_storage_full[511:480];
assign main_genericstandalone_csrbank0_o_data14_w = main_rtio_o_data_storage_full[479:448];
assign main_genericstandalone_csrbank0_o_data13_w = main_rtio_o_data_storage_full[447:416];
assign main_genericstandalone_csrbank0_o_data12_w = main_rtio_o_data_storage_full[415:384];
assign main_genericstandalone_csrbank0_o_data11_w = main_rtio_o_data_storage_full[383:352];
assign main_genericstandalone_csrbank0_o_data10_w = main_rtio_o_data_storage_full[351:320];
assign main_genericstandalone_csrbank0_o_data9_w = main_rtio_o_data_storage_full[319:288];
assign main_genericstandalone_csrbank0_o_data8_w = main_rtio_o_data_storage_full[287:256];
assign main_genericstandalone_csrbank0_o_data7_w = main_rtio_o_data_storage_full[255:224];
assign main_genericstandalone_csrbank0_o_data6_w = main_rtio_o_data_storage_full[223:192];
assign main_genericstandalone_csrbank0_o_data5_w = main_rtio_o_data_storage_full[191:160];
assign main_genericstandalone_csrbank0_o_data4_w = main_rtio_o_data_storage_full[159:128];
assign main_genericstandalone_csrbank0_o_data3_w = main_rtio_o_data_storage_full[127:96];
assign main_genericstandalone_csrbank0_o_data2_w = main_rtio_o_data_storage_full[95:64];
assign main_genericstandalone_csrbank0_o_data1_w = main_rtio_o_data_storage_full[63:32];
assign main_genericstandalone_csrbank0_o_data0_w = main_rtio_o_data_storage_full[31:0];
assign main_genericstandalone_csrbank0_o_status_w = main_rtio_o_status_status[2:0];
assign main_rtio_i_timeout_storage = main_rtio_i_timeout_storage_full[63:0];
assign main_genericstandalone_csrbank0_i_timeout1_w = main_rtio_i_timeout_storage_full[63:32];
assign main_genericstandalone_csrbank0_i_timeout0_w = main_rtio_i_timeout_storage_full[31:0];
assign main_genericstandalone_csrbank0_i_data_w = main_rtio_i_data_status[31:0];
assign main_genericstandalone_csrbank0_i_timestamp1_w = main_rtio_i_timestamp_status[63:32];
assign main_genericstandalone_csrbank0_i_timestamp0_w = main_rtio_i_timestamp_status[31:0];
assign main_genericstandalone_csrbank0_i_status_w = main_rtio_i_status_status[3:0];
assign main_genericstandalone_csrbank0_counter1_w = main_rtio_counter_status[63:32];
assign main_genericstandalone_csrbank0_counter0_w = main_rtio_counter_status[31:0];
assign main_dma_enable_enable_r = main_genericstandalone_csrbank1_bus_dat_w[0];
assign main_dma_enable_enable_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 1'd0));
assign main_genericstandalone_csrbank1_base_address1_r = main_genericstandalone_csrbank1_bus_dat_w[1:0];
assign main_genericstandalone_csrbank1_base_address1_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 1'd1));
assign main_genericstandalone_csrbank1_base_address0_r = main_genericstandalone_csrbank1_bus_dat_w[31:0];
assign main_genericstandalone_csrbank1_base_address0_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 2'd2));
assign main_genericstandalone_csrbank1_time_offset1_r = main_genericstandalone_csrbank1_bus_dat_w[31:0];
assign main_genericstandalone_csrbank1_time_offset1_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 2'd3));
assign main_genericstandalone_csrbank1_time_offset0_r = main_genericstandalone_csrbank1_bus_dat_w[31:0];
assign main_genericstandalone_csrbank1_time_offset0_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 3'd4));
assign main_dma_cri_master_error_r = main_genericstandalone_csrbank1_bus_dat_w[1:0];
assign main_dma_cri_master_error_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 3'd5));
assign main_genericstandalone_csrbank1_error_channel_r = main_genericstandalone_csrbank1_bus_dat_w[23:0];
assign main_genericstandalone_csrbank1_error_channel_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 3'd6));
assign main_genericstandalone_csrbank1_error_timestamp1_r = main_genericstandalone_csrbank1_bus_dat_w[31:0];
assign main_genericstandalone_csrbank1_error_timestamp1_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 3'd7));
assign main_genericstandalone_csrbank1_error_timestamp0_r = main_genericstandalone_csrbank1_bus_dat_w[31:0];
assign main_genericstandalone_csrbank1_error_timestamp0_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 4'd8));
assign main_genericstandalone_csrbank1_error_address_r = main_genericstandalone_csrbank1_bus_dat_w[15:0];
assign main_genericstandalone_csrbank1_error_address_re = ((((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb) & (~main_genericstandalone_csrbank1_bus_ack)) & main_genericstandalone_csrbank1_bus_we) & (main_genericstandalone_csrbank1_bus_adr[3:0] == 4'd9));
assign main_dma_dma_storage = main_dma_dma_storage_full[33:4];
assign main_genericstandalone_csrbank1_base_address1_w = main_dma_dma_storage_full[33:32];
assign main_genericstandalone_csrbank1_base_address0_w = {main_dma_dma_storage_full[31:4], {28{1'd0}}};
assign main_dma_time_offset_storage = main_dma_time_offset_storage_full[63:0];
assign main_genericstandalone_csrbank1_time_offset1_w = main_dma_time_offset_storage_full[63:32];
assign main_genericstandalone_csrbank1_time_offset0_w = main_dma_time_offset_storage_full[31:0];
assign main_genericstandalone_csrbank1_error_channel_w = main_dma_cri_master_error_channel_status[23:0];
assign main_genericstandalone_csrbank1_error_timestamp1_w = main_dma_cri_master_error_timestamp_status[63:32];
assign main_genericstandalone_csrbank1_error_timestamp0_w = main_dma_cri_master_error_timestamp_status[31:0];
assign main_genericstandalone_csrbank1_error_address_w = main_dma_cri_master_error_address_status[15:0];
assign main_cri_con_shared_cmd = builder_comb_rhs_array_muxed10;
assign main_cri_con_shared_chan_sel = builder_comb_rhs_array_muxed11;
assign main_cri_con_shared_o_timestamp = builder_comb_rhs_array_muxed12;
assign main_cri_con_shared_o_data = builder_comb_rhs_array_muxed13;
assign main_cri_con_shared_o_address = builder_comb_rhs_array_muxed14;
assign main_cri_con_shared_i_timeout = builder_comb_rhs_array_muxed15;
assign main_rtio_cri_o_status = main_cri_con_shared_o_status;
assign main_dma_cri_master_cri_o_status = main_cri_con_shared_o_status;
assign main_rtio_cri_o_buffer_space_valid = main_cri_con_shared_o_buffer_space_valid;
assign main_dma_cri_master_cri_o_buffer_space_valid = main_cri_con_shared_o_buffer_space_valid;
assign main_rtio_cri_o_buffer_space = main_cri_con_shared_o_buffer_space;
assign main_dma_cri_master_cri_o_buffer_space = main_cri_con_shared_o_buffer_space;
assign main_rtio_cri_i_data = main_cri_con_shared_i_data;
assign main_dma_cri_master_cri_i_data = main_cri_con_shared_i_data;
assign main_rtio_cri_i_timestamp = main_cri_con_shared_i_timestamp;
assign main_dma_cri_master_cri_i_timestamp = main_cri_con_shared_i_timestamp;
assign main_rtio_cri_i_status = main_cri_con_shared_i_status;
assign main_dma_cri_master_cri_i_status = main_cri_con_shared_i_status;
assign main_rtio_core_cri_chan_sel = main_cri_con_shared_chan_sel;
assign main_rtio_core_cri_o_timestamp = main_cri_con_shared_o_timestamp;
assign main_rtio_core_cri_o_data = main_cri_con_shared_o_data;
assign main_rtio_core_cri_o_address = main_cri_con_shared_o_address;
assign main_rtio_core_cri_i_timeout = main_cri_con_shared_i_timeout;

// synthesis translate_off
reg dummy_d_160;
// synthesis translate_on
always @(*) begin
	main_rtio_core_cri_cmd <= 2'd0;
	if ((main_cri_con_selected == 1'd0)) begin
		main_rtio_core_cri_cmd <= main_cri_con_shared_cmd;
	end
// synthesis translate_off
	dummy_d_160 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_161;
// synthesis translate_on
always @(*) begin
	main_cri_con_shared_o_status <= 3'd0;
	main_cri_con_shared_o_buffer_space_valid <= 1'd0;
	main_cri_con_shared_o_buffer_space <= 16'd0;
	main_cri_con_shared_i_data <= 32'd0;
	main_cri_con_shared_i_timestamp <= 64'd0;
	main_cri_con_shared_i_status <= 4'd0;
	case (main_cri_con_selected)
		1'd0: begin
			main_cri_con_shared_o_status <= main_rtio_core_cri_o_status;
			main_cri_con_shared_o_buffer_space_valid <= main_rtio_core_cri_o_buffer_space_valid;
			main_cri_con_shared_o_buffer_space <= main_rtio_core_cri_o_buffer_space;
			main_cri_con_shared_i_data <= main_rtio_core_cri_i_data;
			main_cri_con_shared_i_timestamp <= main_rtio_core_cri_i_timestamp;
			main_cri_con_shared_i_status <= main_rtio_core_cri_i_status;
		end
	endcase
// synthesis translate_off
	dummy_d_161 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_csrbank2_selected0_r = main_genericstandalone_csrbank2_bus_dat_w[1:0];
assign main_genericstandalone_csrbank2_selected0_re = ((((main_genericstandalone_csrbank2_bus_cyc & main_genericstandalone_csrbank2_bus_stb) & (~main_genericstandalone_csrbank2_bus_ack)) & main_genericstandalone_csrbank2_bus_we) & (main_genericstandalone_csrbank2_bus_adr[0] == 1'd0));
assign main_cri_con_storage = main_cri_con_storage_full[1:0];
assign main_genericstandalone_csrbank2_selected0_w = main_cri_con_storage_full[1:0];
assign main_mon_bussynchronizer0_i = main_inout_8x0_serdes_i0[7];
assign main_mon_bussynchronizer1_i = main_inout_8x0_serdes_oe;
assign main_mon_bussynchronizer2_i = main_inout_8x1_serdes_i0[7];
assign main_mon_bussynchronizer3_i = main_inout_8x1_serdes_oe;
assign main_mon_bussynchronizer4_i = main_inout_8x2_serdes_i0[7];
assign main_mon_bussynchronizer5_i = main_inout_8x2_serdes_oe;
assign main_mon_bussynchronizer6_i = main_inout_8x3_serdes_i0[7];
assign main_mon_bussynchronizer7_i = main_inout_8x3_serdes_oe;
assign main_mon_bussynchronizer8_i = main_inout_8x4_serdes_i0[7];
assign main_mon_bussynchronizer9_i = main_inout_8x4_serdes_oe;
assign main_mon_bussynchronizer10_i = main_inout_8x5_serdes_i0[7];
assign main_mon_bussynchronizer11_i = main_inout_8x5_serdes_oe;
assign main_mon_bussynchronizer12_i = main_inout_8x6_serdes_i0[7];
assign main_mon_bussynchronizer13_i = main_inout_8x6_serdes_oe;
assign main_mon_bussynchronizer14_i = main_inout_8x7_serdes_i0[7];
assign main_mon_bussynchronizer15_i = main_inout_8x7_serdes_oe;
assign main_mon_bussynchronizer16_i = main_output_8x0_o[7];
assign main_mon_bussynchronizer17_i = main_output_8x1_o[7];
assign main_mon_bussynchronizer18_i = main_output_8x2_o[7];
assign main_mon_bussynchronizer19_i = main_output_8x3_o[7];
assign main_mon_bussynchronizer20_i = main_output_8x4_o[7];
assign main_mon_bussynchronizer21_i = main_output_8x5_o[7];
assign main_mon_bussynchronizer22_i = main_output_8x6_o[7];
assign main_mon_bussynchronizer23_i = main_output_8x7_o[7];
assign main_mon_bussynchronizer24_i = main_output_8x8_o[7];
assign main_mon_bussynchronizer25_i = main_output_8x9_o[7];
assign main_mon_bussynchronizer26_i = main_output_8x10_o[7];
assign main_mon_bussynchronizer27_i = main_output_8x11_o[7];
assign main_mon_bussynchronizer28_i = main_output_8x12_o[7];
assign main_mon_bussynchronizer29_i = main_output_8x13_o[7];
assign main_mon_bussynchronizer30_i = main_output_8x14_o[7];
assign main_mon_bussynchronizer31_i = main_output_8x15_o[7];
assign main_mon_bussynchronizer32_i = main_output_8x16_o[7];
assign main_mon_bussynchronizer33_i = main_output_8x17_o[7];
assign main_mon_bussynchronizer34_i = main_output_8x18_o[7];
assign main_mon_bussynchronizer35_i = main_output_8x19_o[7];
assign main_mon_bussynchronizer36_i = main_output_8x20_o[7];
assign main_mon_bussynchronizer37_i = main_output_8x21_o[7];
assign main_mon_bussynchronizer38_i = main_output_8x22_o[7];
assign main_mon_bussynchronizer39_i = main_output0_pad_o;
assign main_mon_bussynchronizer40_i = main_output1_pad_o;
assign main_inj_value_w = builder_comb_rhs_array_muxed16;
assign main_rtio_analyzer_fifo_sink_stb = main_rtio_analyzer_message_encoder_source_stb;
assign main_rtio_analyzer_message_encoder_source_ack = main_rtio_analyzer_fifo_sink_ack;
assign main_rtio_analyzer_fifo_sink_eop = main_rtio_analyzer_message_encoder_source_eop;
assign main_rtio_analyzer_fifo_sink_payload_data = main_rtio_analyzer_message_encoder_source_payload_data;
assign main_rtio_analyzer_converter_sink_stb = main_rtio_analyzer_fifo_source_stb;
assign main_rtio_analyzer_fifo_source_ack = main_rtio_analyzer_converter_sink_ack;
assign main_rtio_analyzer_converter_sink_eop = main_rtio_analyzer_fifo_source_eop;
assign main_rtio_analyzer_converter_sink_payload_data = main_rtio_analyzer_fifo_source_payload_data;
assign main_rtio_analyzer_dma_sink_stb = main_rtio_analyzer_converter_source_stb;
assign main_rtio_analyzer_converter_source_ack = main_rtio_analyzer_dma_sink_ack;
assign main_rtio_analyzer_dma_sink_eop = main_rtio_analyzer_converter_source_eop;
assign main_rtio_analyzer_dma_sink_payload_data = main_rtio_analyzer_converter_source_payload_data;
assign main_rtio_analyzer_dma_sink_payload_valid_token_count = main_rtio_analyzer_converter_source_payload_valid_token_count;

// synthesis translate_off
reg dummy_d_162;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_read_done <= 1'd0;
	main_rtio_analyzer_message_encoder_read_overflow <= 1'd0;
	if ((main_rtio_analyzer_message_encoder_read_wait_event_r & (~main_rtio_core_cri_i_status[2]))) begin
		if ((~main_rtio_core_cri_i_status[0])) begin
			main_rtio_analyzer_message_encoder_read_done <= 1'd1;
		end
		if (main_rtio_core_cri_i_status[1]) begin
			main_rtio_analyzer_message_encoder_read_overflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_162 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_input_output_channel = main_rtio_core_cri_chan_sel;
assign main_rtio_analyzer_message_encoder_input_output_address_padding = main_rtio_core_cri_o_address;
assign main_rtio_analyzer_message_encoder_input_output_rtio_counter = main_rtio_tsc_full_ts_sys;

// synthesis translate_off
reg dummy_d_163;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_input_output_message_type <= 2'd0;
	main_rtio_analyzer_message_encoder_input_output_timestamp <= 64'd0;
	main_rtio_analyzer_message_encoder_input_output_data <= 64'd0;
	if ((main_rtio_core_cri_cmd == 1'd1)) begin
		main_rtio_analyzer_message_encoder_input_output_message_type <= 1'd0;
		main_rtio_analyzer_message_encoder_input_output_timestamp <= main_rtio_core_cri_o_timestamp;
		main_rtio_analyzer_message_encoder_input_output_data <= main_rtio_core_cri_o_data;
	end else begin
		main_rtio_analyzer_message_encoder_input_output_message_type <= 1'd1;
		main_rtio_analyzer_message_encoder_input_output_timestamp <= main_rtio_core_cri_i_timestamp;
		main_rtio_analyzer_message_encoder_input_output_data <= main_rtio_core_cri_i_data;
	end
// synthesis translate_off
	dummy_d_163 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_input_output_stb = ((main_rtio_core_cri_cmd == 1'd1) | main_rtio_analyzer_message_encoder_read_done);
assign main_rtio_analyzer_message_encoder_exception_message_type = 2'd2;
assign main_rtio_analyzer_message_encoder_exception_channel = main_rtio_core_cri_chan_sel;
assign main_rtio_analyzer_message_encoder_exception_rtio_counter = main_rtio_tsc_full_ts_sys;

// synthesis translate_off
reg dummy_d_164;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_exception_stb <= 1'd0;
	main_rtio_analyzer_message_encoder_exception_exception_type <= 8'd0;
	if ((main_rtio_analyzer_message_encoder_just_written & main_rtio_core_cri_o_status[1])) begin
		main_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_rtio_analyzer_message_encoder_exception_exception_type <= 5'd20;
	end
	if (main_rtio_analyzer_message_encoder_read_overflow) begin
		main_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_rtio_analyzer_message_encoder_exception_exception_type <= 6'd33;
	end
// synthesis translate_off
	dummy_d_164 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_stopped_message_type = 2'd3;
assign main_rtio_analyzer_message_encoder_stopped_rtio_counter = main_rtio_tsc_full_ts_sys;
assign main_rtio_analyzer_fifo_syncfifo_din = {main_rtio_analyzer_fifo_fifo_in_eop, main_rtio_analyzer_fifo_fifo_in_payload_data};
assign {main_rtio_analyzer_fifo_fifo_out_eop, main_rtio_analyzer_fifo_fifo_out_payload_data} = main_rtio_analyzer_fifo_syncfifo_dout;
assign main_rtio_analyzer_fifo_sink_ack = main_rtio_analyzer_fifo_syncfifo_writable;
assign main_rtio_analyzer_fifo_syncfifo_we = main_rtio_analyzer_fifo_sink_stb;
assign main_rtio_analyzer_fifo_fifo_in_eop = main_rtio_analyzer_fifo_sink_eop;
assign main_rtio_analyzer_fifo_fifo_in_payload_data = main_rtio_analyzer_fifo_sink_payload_data;
assign main_rtio_analyzer_fifo_source_stb = main_rtio_analyzer_fifo_readable;
assign main_rtio_analyzer_fifo_source_eop = main_rtio_analyzer_fifo_fifo_out_eop;
assign main_rtio_analyzer_fifo_source_payload_data = main_rtio_analyzer_fifo_fifo_out_payload_data;
assign main_rtio_analyzer_fifo_re = main_rtio_analyzer_fifo_source_ack;
assign main_rtio_analyzer_fifo_syncfifo_re = (main_rtio_analyzer_fifo_syncfifo_readable & ((~main_rtio_analyzer_fifo_readable) | main_rtio_analyzer_fifo_re));
assign main_rtio_analyzer_fifo_level1 = (main_rtio_analyzer_fifo_level0 + main_rtio_analyzer_fifo_readable);

// synthesis translate_off
reg dummy_d_165;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_fifo_wrport_adr <= 7'd0;
	if (main_rtio_analyzer_fifo_replace) begin
		main_rtio_analyzer_fifo_wrport_adr <= (main_rtio_analyzer_fifo_produce - 1'd1);
	end else begin
		main_rtio_analyzer_fifo_wrport_adr <= main_rtio_analyzer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_165 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_fifo_wrport_dat_w = main_rtio_analyzer_fifo_syncfifo_din;
assign main_rtio_analyzer_fifo_wrport_we = (main_rtio_analyzer_fifo_syncfifo_we & (main_rtio_analyzer_fifo_syncfifo_writable | main_rtio_analyzer_fifo_replace));
assign main_rtio_analyzer_fifo_do_read = (main_rtio_analyzer_fifo_syncfifo_readable & main_rtio_analyzer_fifo_syncfifo_re);
assign main_rtio_analyzer_fifo_rdport_adr = main_rtio_analyzer_fifo_consume;
assign main_rtio_analyzer_fifo_syncfifo_dout = main_rtio_analyzer_fifo_rdport_dat_r;
assign main_rtio_analyzer_fifo_rdport_re = main_rtio_analyzer_fifo_do_read;
assign main_rtio_analyzer_fifo_syncfifo_writable = (main_rtio_analyzer_fifo_level0 != 8'd128);
assign main_rtio_analyzer_fifo_syncfifo_readable = (main_rtio_analyzer_fifo_level0 != 1'd0);
assign main_rtio_analyzer_converter_last = (main_rtio_analyzer_converter_mux == 1'd1);
assign main_rtio_analyzer_converter_source_stb = main_rtio_analyzer_converter_sink_stb;
assign main_rtio_analyzer_converter_source_eop = (main_rtio_analyzer_converter_sink_eop & main_rtio_analyzer_converter_last);
assign main_rtio_analyzer_converter_sink_ack = (main_rtio_analyzer_converter_last & main_rtio_analyzer_converter_source_ack);

// synthesis translate_off
reg dummy_d_166;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_converter_source_payload_data <= 128'd0;
	case (main_rtio_analyzer_converter_mux)
		1'd0: begin
			main_rtio_analyzer_converter_source_payload_data <= main_rtio_analyzer_converter_sink_payload_data[255:128];
		end
		default: begin
			main_rtio_analyzer_converter_source_payload_data <= main_rtio_analyzer_converter_sink_payload_data[127:0];
		end
	endcase
// synthesis translate_off
	dummy_d_166 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_converter_source_payload_valid_token_count = main_rtio_analyzer_converter_last;
assign main_genericstandalone_interface1_bus_cyc = main_rtio_analyzer_dma_sink_stb;
assign main_genericstandalone_interface1_bus_stb = main_rtio_analyzer_dma_sink_stb;
assign main_rtio_analyzer_dma_sink_ack = main_genericstandalone_interface1_bus_ack;
assign main_genericstandalone_interface1_bus_we = 1'd1;
assign main_genericstandalone_interface1_bus_dat_w = main_rtio_analyzer_dma_sink_payload_data;
assign main_genericstandalone_interface1_bus_sel = 16'd65535;
assign main_rtio_analyzer_dma_status = (main_rtio_analyzer_dma_message_count <<< 3'd5);
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr = builder_comb_rhs_array_muxed54;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_w = builder_comb_rhs_array_muxed55;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_sel = builder_comb_rhs_array_muxed56;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cyc = builder_comb_rhs_array_muxed57;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_stb = builder_comb_rhs_array_muxed58;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_we = builder_comb_rhs_array_muxed59;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_cti = builder_comb_rhs_array_muxed60;
assign main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_bte = builder_comb_rhs_array_muxed61;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
assign main_genericstandalone_kernel_cpu_wb_sdram_dat_r = main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_wb_sdram_ack = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_genericstandalone_kernel_cpu_wb_sdram_err = (main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign builder_sdram_cpulevel_arbiter_request = {(main_genericstandalone_kernel_cpu_wb_sdram_cyc & (~main_genericstandalone_kernel_cpu_wb_sdram_ack)), (main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc & (~main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack))};
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_adr = builder_comb_rhs_array_muxed62;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_w = builder_comb_rhs_array_muxed63;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_sel = builder_comb_rhs_array_muxed64;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cyc = builder_comb_rhs_array_muxed65;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_stb = builder_comb_rhs_array_muxed66;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_we = builder_comb_rhs_array_muxed67;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_cti = builder_comb_rhs_array_muxed68;
assign main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_bte = builder_comb_rhs_array_muxed69;
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_interface0_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_interface1_bus_dat_r = main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_genericstandalone_interface0_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_genericstandalone_interface1_bus_ack = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 2'd2));
assign main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_genericstandalone_interface0_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_genericstandalone_interface1_bus_err = (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 2'd2));
assign builder_sdram_native_arbiter_request = {(main_genericstandalone_interface1_bus_cyc & (~main_genericstandalone_interface1_bus_ack)), (main_genericstandalone_interface0_bus_cyc & (~main_genericstandalone_interface0_bus_ack)), (main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc & (~main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_ack))};
assign builder_genericstandalone_shared_adr = builder_comb_rhs_array_muxed70;
assign builder_genericstandalone_shared_dat_w = builder_comb_rhs_array_muxed71;
assign builder_genericstandalone_shared_sel = builder_comb_rhs_array_muxed72;
assign builder_genericstandalone_shared_cyc = builder_comb_rhs_array_muxed73;
assign builder_genericstandalone_shared_stb = builder_comb_rhs_array_muxed74;
assign builder_genericstandalone_shared_we = builder_comb_rhs_array_muxed75;
assign builder_genericstandalone_shared_cti = builder_comb_rhs_array_muxed76;
assign builder_genericstandalone_shared_bte = builder_comb_rhs_array_muxed77;
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r = builder_genericstandalone_shared_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_r = builder_genericstandalone_shared_dat_r;
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_ack = (builder_genericstandalone_shared_ack & (builder_genericstandalone_grant == 1'd0));
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_ack = (builder_genericstandalone_shared_ack & (builder_genericstandalone_grant == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_ibus_err = (builder_genericstandalone_shared_err & (builder_genericstandalone_grant == 1'd0));
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_err = (builder_genericstandalone_shared_err & (builder_genericstandalone_grant == 1'd1));
assign builder_genericstandalone_request = {(main_genericstandalone_genericstandalone_genericstandalone_tmpu_cyc & (~main_genericstandalone_genericstandalone_genericstandalone_tmpu_ack)), (main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc & (~main_genericstandalone_genericstandalone_genericstandalone_ibus_ack))};

// synthesis translate_off
reg dummy_d_167;
// synthesis translate_on
always @(*) begin
	builder_genericstandalone_slave_sel <= 6'd0;
	builder_genericstandalone_slave_sel[0] <= (((1'd1 & (~builder_genericstandalone_shared_adr[27])) & (~builder_genericstandalone_shared_adr[28])) & builder_genericstandalone_shared_adr[26]);
	builder_genericstandalone_slave_sel[1] <= (((1'd1 & (~builder_genericstandalone_shared_adr[26])) & builder_genericstandalone_shared_adr[27]) & builder_genericstandalone_shared_adr[28]);
	builder_genericstandalone_slave_sel[2] <= ((1'd1 & (~builder_genericstandalone_shared_adr[27])) & builder_genericstandalone_shared_adr[28]);
	builder_genericstandalone_slave_sel[3] <= (((1'd1 & (~builder_genericstandalone_shared_adr[26])) & (~builder_genericstandalone_shared_adr[27])) & (~builder_genericstandalone_shared_adr[28]));
	builder_genericstandalone_slave_sel[4] <= ((1'd1 & (~builder_genericstandalone_shared_adr[28])) & builder_genericstandalone_shared_adr[27]);
	builder_genericstandalone_slave_sel[5] <= (((1'd1 & builder_genericstandalone_shared_adr[26]) & builder_genericstandalone_shared_adr[27]) & builder_genericstandalone_shared_adr[28]);
// synthesis translate_off
	dummy_d_167 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_spiflash_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_genericstandalone_spiflash_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_genericstandalone_spiflash_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_genericstandalone_spiflash_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_genericstandalone_spiflash_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_genericstandalone_spiflash_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_genericstandalone_spiflash_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_bus_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_bus_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_bus_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_bus_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_bus_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_bus_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_bus_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_mailbox_i1_adr = builder_genericstandalone_shared_adr;
assign main_genericstandalone_mailbox_i1_dat_w = builder_genericstandalone_shared_dat_w;
assign main_genericstandalone_mailbox_i1_sel = builder_genericstandalone_shared_sel;
assign main_genericstandalone_mailbox_i1_stb = builder_genericstandalone_shared_stb;
assign main_genericstandalone_mailbox_i1_we = builder_genericstandalone_shared_we;
assign main_genericstandalone_mailbox_i1_cti = builder_genericstandalone_shared_cti;
assign main_genericstandalone_mailbox_i1_bte = builder_genericstandalone_shared_bte;
assign main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[0]);
assign main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[1]);
assign main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[2]);
assign main_genericstandalone_genericstandalone_spiflash_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[3]);
assign main_genericstandalone_bus_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[4]);
assign main_genericstandalone_mailbox_i1_cyc = (builder_genericstandalone_shared_cyc & builder_genericstandalone_slave_sel[5]);
assign builder_genericstandalone_shared_ack = (((((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack | main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack) | main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_ack) | main_genericstandalone_genericstandalone_spiflash_bus_ack) | main_genericstandalone_bus_ack) | main_genericstandalone_mailbox_i1_ack);
assign builder_genericstandalone_shared_err = (((((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_err | main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_err) | main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_err) | main_genericstandalone_genericstandalone_spiflash_bus_err) | main_genericstandalone_bus_err) | main_genericstandalone_mailbox_i1_err);
assign builder_genericstandalone_shared_dat_r = (((((({32{builder_genericstandalone_slave_sel_r[0]}} & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_dat_r) | ({32{builder_genericstandalone_slave_sel_r[1]}} & main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r)) | ({32{builder_genericstandalone_slave_sel_r[2]}} & main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_r)) | ({32{builder_genericstandalone_slave_sel_r[3]}} & main_genericstandalone_genericstandalone_spiflash_bus_dat_r)) | ({32{builder_genericstandalone_slave_sel_r[4]}} & main_genericstandalone_bus_dat_r)) | ({32{builder_genericstandalone_slave_sel_r[5]}} & main_genericstandalone_mailbox_i1_dat_r));
assign builder_genericstandalone_csrbank0_sel = (builder_genericstandalone_interface0_bank_bus_adr[13:9] == 3'd7);
assign builder_genericstandalone_csrbank0_dly_sel0_r = builder_genericstandalone_interface0_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank0_dly_sel0_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[1:0] == 1'd0));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_r = builder_genericstandalone_interface0_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[1:0] == 1'd1));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_r = builder_genericstandalone_interface0_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[1:0] == 2'd2));
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_r = builder_genericstandalone_interface0_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re = ((builder_genericstandalone_csrbank0_sel & builder_genericstandalone_interface0_bank_bus_we) & (builder_genericstandalone_interface0_bank_bus_adr[1:0] == 2'd3));
assign main_genericstandalone_genericstandalone_ddrphy_storage = main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0];
assign builder_genericstandalone_csrbank0_dly_sel0_w = main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0];
assign builder_genericstandalone_csrbank1_sel = (builder_genericstandalone_interface1_bank_bus_adr[13:9] == 3'd5);
assign builder_genericstandalone_csrbank1_control0_r = builder_genericstandalone_interface1_bank_bus_dat_w[3:0];
assign builder_genericstandalone_csrbank1_control0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 1'd0));
assign builder_genericstandalone_csrbank1_pi0_command0_r = builder_genericstandalone_interface1_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank1_pi0_command0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 1'd1));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 2'd2));
assign builder_genericstandalone_csrbank1_pi0_address1_r = builder_genericstandalone_interface1_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank1_pi0_address1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 2'd3));
assign builder_genericstandalone_csrbank1_pi0_address0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_address0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 3'd4));
assign builder_genericstandalone_csrbank1_pi0_baddress0_r = builder_genericstandalone_interface1_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank1_pi0_baddress0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 3'd5));
assign builder_genericstandalone_csrbank1_pi0_wrdata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_wrdata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 3'd6));
assign builder_genericstandalone_csrbank1_pi0_wrdata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_wrdata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 3'd7));
assign builder_genericstandalone_csrbank1_pi0_wrdata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_wrdata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd8));
assign builder_genericstandalone_csrbank1_pi0_wrdata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_wrdata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd9));
assign builder_genericstandalone_csrbank1_pi0_rddata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_rddata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd10));
assign builder_genericstandalone_csrbank1_pi0_rddata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_rddata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd11));
assign builder_genericstandalone_csrbank1_pi0_rddata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_rddata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd12));
assign builder_genericstandalone_csrbank1_pi0_rddata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi0_rddata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd13));
assign builder_genericstandalone_csrbank1_pi1_command0_r = builder_genericstandalone_interface1_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank1_pi1_command0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd14));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 4'd15));
assign builder_genericstandalone_csrbank1_pi1_address1_r = builder_genericstandalone_interface1_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank1_pi1_address1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd16));
assign builder_genericstandalone_csrbank1_pi1_address0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_address0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd17));
assign builder_genericstandalone_csrbank1_pi1_baddress0_r = builder_genericstandalone_interface1_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank1_pi1_baddress0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd18));
assign builder_genericstandalone_csrbank1_pi1_wrdata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_wrdata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd19));
assign builder_genericstandalone_csrbank1_pi1_wrdata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_wrdata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd20));
assign builder_genericstandalone_csrbank1_pi1_wrdata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_wrdata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd21));
assign builder_genericstandalone_csrbank1_pi1_wrdata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_wrdata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd22));
assign builder_genericstandalone_csrbank1_pi1_rddata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_rddata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd23));
assign builder_genericstandalone_csrbank1_pi1_rddata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_rddata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd24));
assign builder_genericstandalone_csrbank1_pi1_rddata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_rddata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd25));
assign builder_genericstandalone_csrbank1_pi1_rddata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi1_rddata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd26));
assign builder_genericstandalone_csrbank1_pi2_command0_r = builder_genericstandalone_interface1_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank1_pi2_command0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd27));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd28));
assign builder_genericstandalone_csrbank1_pi2_address1_r = builder_genericstandalone_interface1_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank1_pi2_address1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd29));
assign builder_genericstandalone_csrbank1_pi2_address0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_address0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd30));
assign builder_genericstandalone_csrbank1_pi2_baddress0_r = builder_genericstandalone_interface1_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank1_pi2_baddress0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 5'd31));
assign builder_genericstandalone_csrbank1_pi2_wrdata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_wrdata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd32));
assign builder_genericstandalone_csrbank1_pi2_wrdata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_wrdata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd33));
assign builder_genericstandalone_csrbank1_pi2_wrdata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_wrdata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd34));
assign builder_genericstandalone_csrbank1_pi2_wrdata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_wrdata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd35));
assign builder_genericstandalone_csrbank1_pi2_rddata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_rddata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd36));
assign builder_genericstandalone_csrbank1_pi2_rddata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_rddata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd37));
assign builder_genericstandalone_csrbank1_pi2_rddata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_rddata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd38));
assign builder_genericstandalone_csrbank1_pi2_rddata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi2_rddata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd39));
assign builder_genericstandalone_csrbank1_pi3_command0_r = builder_genericstandalone_interface1_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank1_pi3_command0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd40));
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_r = builder_genericstandalone_interface1_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd41));
assign builder_genericstandalone_csrbank1_pi3_address1_r = builder_genericstandalone_interface1_bank_bus_dat_w[6:0];
assign builder_genericstandalone_csrbank1_pi3_address1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd42));
assign builder_genericstandalone_csrbank1_pi3_address0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_address0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd43));
assign builder_genericstandalone_csrbank1_pi3_baddress0_r = builder_genericstandalone_interface1_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank1_pi3_baddress0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd44));
assign builder_genericstandalone_csrbank1_pi3_wrdata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_wrdata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd45));
assign builder_genericstandalone_csrbank1_pi3_wrdata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_wrdata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd46));
assign builder_genericstandalone_csrbank1_pi3_wrdata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_wrdata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd47));
assign builder_genericstandalone_csrbank1_pi3_wrdata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_wrdata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd48));
assign builder_genericstandalone_csrbank1_pi3_rddata3_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_rddata3_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd49));
assign builder_genericstandalone_csrbank1_pi3_rddata2_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_rddata2_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd50));
assign builder_genericstandalone_csrbank1_pi3_rddata1_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_rddata1_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd51));
assign builder_genericstandalone_csrbank1_pi3_rddata0_r = builder_genericstandalone_interface1_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank1_pi3_rddata0_re = ((builder_genericstandalone_csrbank1_sel & builder_genericstandalone_interface1_bank_bus_we) & (builder_genericstandalone_interface1_bank_bus_adr[5:0] == 6'd52));
assign main_genericstandalone_genericstandalone_genericstandalone_storage = main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0];
assign builder_genericstandalone_csrbank1_control0_w = main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0];
assign builder_genericstandalone_csrbank1_pi0_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:0];
assign builder_genericstandalone_csrbank1_pi0_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:8];
assign builder_genericstandalone_csrbank1_pi0_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank1_pi0_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank1_pi0_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank1_pi0_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank1_pi0_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank1_pi0_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank1_pi0_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[31:24];
assign builder_genericstandalone_csrbank1_pi0_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[23:16];
assign builder_genericstandalone_csrbank1_pi0_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[15:8];
assign builder_genericstandalone_csrbank1_pi0_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0];
assign builder_genericstandalone_csrbank1_pi1_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:0];
assign builder_genericstandalone_csrbank1_pi1_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:8];
assign builder_genericstandalone_csrbank1_pi1_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank1_pi1_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank1_pi1_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank1_pi1_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank1_pi1_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank1_pi1_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank1_pi1_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[31:24];
assign builder_genericstandalone_csrbank1_pi1_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[23:16];
assign builder_genericstandalone_csrbank1_pi1_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[15:8];
assign builder_genericstandalone_csrbank1_pi1_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0];
assign builder_genericstandalone_csrbank1_pi2_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:0];
assign builder_genericstandalone_csrbank1_pi2_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:8];
assign builder_genericstandalone_csrbank1_pi2_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank1_pi2_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank1_pi2_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank1_pi2_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank1_pi2_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank1_pi2_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank1_pi2_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[31:24];
assign builder_genericstandalone_csrbank1_pi2_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[23:16];
assign builder_genericstandalone_csrbank1_pi2_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[15:8];
assign builder_genericstandalone_csrbank1_pi2_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0];
assign builder_genericstandalone_csrbank1_pi3_command0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:0];
assign builder_genericstandalone_csrbank1_pi3_address1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:8];
assign builder_genericstandalone_csrbank1_pi3_address0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0];
assign builder_genericstandalone_csrbank1_pi3_baddress0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0];
assign main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:0];
assign builder_genericstandalone_csrbank1_pi3_wrdata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:24];
assign builder_genericstandalone_csrbank1_pi3_wrdata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[23:16];
assign builder_genericstandalone_csrbank1_pi3_wrdata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[15:8];
assign builder_genericstandalone_csrbank1_pi3_wrdata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[7:0];
assign builder_genericstandalone_csrbank1_pi3_rddata3_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[31:24];
assign builder_genericstandalone_csrbank1_pi3_rddata2_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[23:16];
assign builder_genericstandalone_csrbank1_pi3_rddata1_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[15:8];
assign builder_genericstandalone_csrbank1_pi3_rddata0_w = main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status[7:0];
assign builder_genericstandalone_csrbank2_sel = (builder_genericstandalone_interface2_bank_bus_adr[13:9] == 4'd10);
assign builder_genericstandalone_csrbank2_sram_writer_slot_r = builder_genericstandalone_interface2_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank2_sram_writer_slot_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank2_sram_writer_length3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_length3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank2_sram_writer_length2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_length2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 2'd2));
assign builder_genericstandalone_csrbank2_sram_writer_length1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_length1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 2'd3));
assign builder_genericstandalone_csrbank2_sram_writer_length0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_length0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank2_sram_writer_errors3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_errors3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank2_sram_writer_errors2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_errors2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 3'd6));
assign builder_genericstandalone_csrbank2_sram_writer_errors1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_errors1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 3'd7));
assign builder_genericstandalone_csrbank2_sram_writer_errors0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_errors0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd8));
assign main_genericstandalone_writer_status_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_writer_status_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd9));
assign main_genericstandalone_writer_pending_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_writer_pending_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank2_sram_writer_ev_enable0_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank2_sram_writer_ev_enable0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd11));
assign main_genericstandalone_reader_start_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_reader_start_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank2_sram_reader_ready_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank2_sram_reader_ready_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank2_sram_reader_slot0_r = builder_genericstandalone_interface2_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank2_sram_reader_slot0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd14));
assign builder_genericstandalone_csrbank2_sram_reader_length1_r = builder_genericstandalone_interface2_bank_bus_dat_w[2:0];
assign builder_genericstandalone_csrbank2_sram_reader_length1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 4'd15));
assign builder_genericstandalone_csrbank2_sram_reader_length0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_sram_reader_length0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd16));
assign main_genericstandalone_reader_eventmanager_status_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_reader_eventmanager_status_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd17));
assign main_genericstandalone_reader_eventmanager_pending_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign main_genericstandalone_reader_eventmanager_pending_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank2_sram_reader_ev_enable0_r = builder_genericstandalone_interface2_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank2_sram_reader_ev_enable0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank2_preamble_errors3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_preamble_errors3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank2_preamble_errors2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_preamble_errors2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank2_preamble_errors1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_preamble_errors1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd22));
assign builder_genericstandalone_csrbank2_preamble_errors0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_preamble_errors0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd23));
assign builder_genericstandalone_csrbank2_crc_errors3_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_crc_errors3_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd24));
assign builder_genericstandalone_csrbank2_crc_errors2_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_crc_errors2_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd25));
assign builder_genericstandalone_csrbank2_crc_errors1_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_crc_errors1_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd26));
assign builder_genericstandalone_csrbank2_crc_errors0_r = builder_genericstandalone_interface2_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank2_crc_errors0_re = ((builder_genericstandalone_csrbank2_sel & builder_genericstandalone_interface2_bank_bus_we) & (builder_genericstandalone_interface2_bank_bus_adr[4:0] == 5'd27));
assign builder_genericstandalone_csrbank2_sram_writer_slot_w = main_genericstandalone_writer_slot_status[1:0];
assign builder_genericstandalone_csrbank2_sram_writer_length3_w = main_genericstandalone_writer_length_status[31:24];
assign builder_genericstandalone_csrbank2_sram_writer_length2_w = main_genericstandalone_writer_length_status[23:16];
assign builder_genericstandalone_csrbank2_sram_writer_length1_w = main_genericstandalone_writer_length_status[15:8];
assign builder_genericstandalone_csrbank2_sram_writer_length0_w = main_genericstandalone_writer_length_status[7:0];
assign builder_genericstandalone_csrbank2_sram_writer_errors3_w = main_genericstandalone_writer_errors_status[31:24];
assign builder_genericstandalone_csrbank2_sram_writer_errors2_w = main_genericstandalone_writer_errors_status[23:16];
assign builder_genericstandalone_csrbank2_sram_writer_errors1_w = main_genericstandalone_writer_errors_status[15:8];
assign builder_genericstandalone_csrbank2_sram_writer_errors0_w = main_genericstandalone_writer_errors_status[7:0];
assign main_genericstandalone_writer_storage = main_genericstandalone_writer_storage_full;
assign builder_genericstandalone_csrbank2_sram_writer_ev_enable0_w = main_genericstandalone_writer_storage_full;
assign builder_genericstandalone_csrbank2_sram_reader_ready_w = main_genericstandalone_reader_ready_status;
assign main_genericstandalone_reader_slot_storage = main_genericstandalone_reader_slot_storage_full[1:0];
assign builder_genericstandalone_csrbank2_sram_reader_slot0_w = main_genericstandalone_reader_slot_storage_full[1:0];
assign main_genericstandalone_reader_length_storage = main_genericstandalone_reader_length_storage_full[10:0];
assign builder_genericstandalone_csrbank2_sram_reader_length1_w = main_genericstandalone_reader_length_storage_full[10:8];
assign builder_genericstandalone_csrbank2_sram_reader_length0_w = main_genericstandalone_reader_length_storage_full[7:0];
assign main_genericstandalone_reader_eventmanager_storage = main_genericstandalone_reader_eventmanager_storage_full;
assign builder_genericstandalone_csrbank2_sram_reader_ev_enable0_w = main_genericstandalone_reader_eventmanager_storage_full;
assign builder_genericstandalone_csrbank2_preamble_errors3_w = main_genericstandalone_preamble_errors_status[31:24];
assign builder_genericstandalone_csrbank2_preamble_errors2_w = main_genericstandalone_preamble_errors_status[23:16];
assign builder_genericstandalone_csrbank2_preamble_errors1_w = main_genericstandalone_preamble_errors_status[15:8];
assign builder_genericstandalone_csrbank2_preamble_errors0_w = main_genericstandalone_preamble_errors_status[7:0];
assign builder_genericstandalone_csrbank2_crc_errors3_w = main_genericstandalone_crc_errors_status[31:24];
assign builder_genericstandalone_csrbank2_crc_errors2_w = main_genericstandalone_crc_errors_status[23:16];
assign builder_genericstandalone_csrbank2_crc_errors1_w = main_genericstandalone_crc_errors_status[15:8];
assign builder_genericstandalone_csrbank2_crc_errors0_w = main_genericstandalone_crc_errors_status[7:0];
assign builder_genericstandalone_csrbank3_sel = (builder_genericstandalone_interface3_bank_bus_adr[13:9] == 4'd13);
assign builder_genericstandalone_csrbank3_in_r = builder_genericstandalone_interface3_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank3_in_re = ((builder_genericstandalone_csrbank3_sel & builder_genericstandalone_interface3_bank_bus_we) & (builder_genericstandalone_interface3_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank3_out0_r = builder_genericstandalone_interface3_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank3_out0_re = ((builder_genericstandalone_csrbank3_sel & builder_genericstandalone_interface3_bank_bus_we) & (builder_genericstandalone_interface3_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank3_oe0_r = builder_genericstandalone_interface3_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank3_oe0_re = ((builder_genericstandalone_csrbank3_sel & builder_genericstandalone_interface3_bank_bus_we) & (builder_genericstandalone_interface3_bank_bus_adr[1:0] == 2'd2));
assign builder_genericstandalone_csrbank3_in_w = main_i2c_status0[1:0];
assign main_i2c_out_storage = main_i2c_out_storage_full[1:0];
assign builder_genericstandalone_csrbank3_out0_w = main_i2c_out_storage_full[1:0];
assign main_i2c_oe_storage = main_i2c_oe_storage_full[1:0];
assign builder_genericstandalone_csrbank3_oe0_w = main_i2c_oe_storage_full[1:0];
assign builder_genericstandalone_csrbank4_sel = (builder_genericstandalone_interface4_bank_bus_adr[13:9] == 2'd2);
assign builder_genericstandalone_csrbank4_address0_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_address0_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank4_data_r = builder_genericstandalone_interface4_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank4_data_re = ((builder_genericstandalone_csrbank4_sel & builder_genericstandalone_interface4_bank_bus_we) & (builder_genericstandalone_interface4_bank_bus_adr[0] == 1'd1));
assign main_add_identifier_storage = main_add_identifier_storage_full[7:0];
assign builder_genericstandalone_csrbank4_address0_w = main_add_identifier_storage_full[7:0];
assign builder_genericstandalone_csrbank4_data_w = main_add_identifier_status[7:0];
assign builder_genericstandalone_csrbank5_sel = (builder_genericstandalone_interface5_bank_bus_adr[13:9] == 4'd11);
assign builder_genericstandalone_csrbank5_reset0_r = builder_genericstandalone_interface5_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank5_reset0_re = ((builder_genericstandalone_csrbank5_sel & builder_genericstandalone_interface5_bank_bus_we) & (builder_genericstandalone_interface5_bank_bus_adr[0] == 1'd0));
assign main_genericstandalone_kernel_cpu_storage = main_genericstandalone_kernel_cpu_storage_full;
assign builder_genericstandalone_csrbank5_reset0_w = main_genericstandalone_kernel_cpu_storage_full;
assign builder_genericstandalone_csrbank6_sel = (builder_genericstandalone_interface6_bank_bus_adr[13:9] == 4'd12);
assign builder_genericstandalone_csrbank6_out0_r = builder_genericstandalone_interface6_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank6_out0_re = ((builder_genericstandalone_csrbank6_sel & builder_genericstandalone_interface6_bank_bus_we) & (builder_genericstandalone_interface6_bank_bus_adr[0] == 1'd0));
assign main_leds_storage = main_leds_storage_full;
assign builder_genericstandalone_csrbank6_out0_w = main_leds_storage_full;
assign builder_genericstandalone_csrbank7_sel = (builder_genericstandalone_interface7_bank_bus_adr[13:9] == 5'd17);
assign builder_genericstandalone_csrbank7_enable0_r = builder_genericstandalone_interface7_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank7_enable0_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank7_busy_r = builder_genericstandalone_interface7_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank7_busy_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank7_message_encoder_overflow_r = builder_genericstandalone_interface7_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank7_message_encoder_overflow_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 2'd2));
assign main_rtio_analyzer_message_encoder_overflow_reset_r = builder_genericstandalone_interface7_bank_bus_dat_w[0];
assign main_rtio_analyzer_message_encoder_overflow_reset_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 2'd3));
assign main_rtio_analyzer_dma_reset_r = builder_genericstandalone_interface7_bank_bus_dat_w[0];
assign main_rtio_analyzer_dma_reset_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank7_dma_base_address4_r = builder_genericstandalone_interface7_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank7_dma_base_address4_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank7_dma_base_address3_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_base_address3_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 3'd6));
assign builder_genericstandalone_csrbank7_dma_base_address2_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_base_address2_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 3'd7));
assign builder_genericstandalone_csrbank7_dma_base_address1_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_base_address1_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd8));
assign builder_genericstandalone_csrbank7_dma_base_address0_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_base_address0_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd9));
assign builder_genericstandalone_csrbank7_dma_last_address4_r = builder_genericstandalone_interface7_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank7_dma_last_address4_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank7_dma_last_address3_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_last_address3_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd11));
assign builder_genericstandalone_csrbank7_dma_last_address2_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_last_address2_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank7_dma_last_address1_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_last_address1_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank7_dma_last_address0_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_last_address0_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd14));
assign builder_genericstandalone_csrbank7_dma_byte_count7_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count7_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 4'd15));
assign builder_genericstandalone_csrbank7_dma_byte_count6_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count6_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd16));
assign builder_genericstandalone_csrbank7_dma_byte_count5_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count5_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd17));
assign builder_genericstandalone_csrbank7_dma_byte_count4_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count4_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank7_dma_byte_count3_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count3_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank7_dma_byte_count2_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count2_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank7_dma_byte_count1_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count1_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank7_dma_byte_count0_r = builder_genericstandalone_interface7_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank7_dma_byte_count0_re = ((builder_genericstandalone_csrbank7_sel & builder_genericstandalone_interface7_bank_bus_we) & (builder_genericstandalone_interface7_bank_bus_adr[4:0] == 5'd22));
assign main_rtio_analyzer_enable_storage = main_rtio_analyzer_enable_storage_full;
assign builder_genericstandalone_csrbank7_enable0_w = main_rtio_analyzer_enable_storage_full;
assign builder_genericstandalone_csrbank7_busy_w = main_rtio_analyzer_busy_status;
assign builder_genericstandalone_csrbank7_message_encoder_overflow_w = main_rtio_analyzer_message_encoder_status;
assign main_rtio_analyzer_dma_base_address_storage = main_rtio_analyzer_dma_base_address_storage_full[33:4];
assign builder_genericstandalone_csrbank7_dma_base_address4_w = main_rtio_analyzer_dma_base_address_storage_full[33:32];
assign builder_genericstandalone_csrbank7_dma_base_address3_w = main_rtio_analyzer_dma_base_address_storage_full[31:24];
assign builder_genericstandalone_csrbank7_dma_base_address2_w = main_rtio_analyzer_dma_base_address_storage_full[23:16];
assign builder_genericstandalone_csrbank7_dma_base_address1_w = main_rtio_analyzer_dma_base_address_storage_full[15:8];
assign builder_genericstandalone_csrbank7_dma_base_address0_w = {main_rtio_analyzer_dma_base_address_storage_full[7:4], {4{1'd0}}};
assign main_rtio_analyzer_dma_last_address_storage = main_rtio_analyzer_dma_last_address_storage_full[33:4];
assign builder_genericstandalone_csrbank7_dma_last_address4_w = main_rtio_analyzer_dma_last_address_storage_full[33:32];
assign builder_genericstandalone_csrbank7_dma_last_address3_w = main_rtio_analyzer_dma_last_address_storage_full[31:24];
assign builder_genericstandalone_csrbank7_dma_last_address2_w = main_rtio_analyzer_dma_last_address_storage_full[23:16];
assign builder_genericstandalone_csrbank7_dma_last_address1_w = main_rtio_analyzer_dma_last_address_storage_full[15:8];
assign builder_genericstandalone_csrbank7_dma_last_address0_w = {main_rtio_analyzer_dma_last_address_storage_full[7:4], {4{1'd0}}};
assign builder_genericstandalone_csrbank7_dma_byte_count7_w = main_rtio_analyzer_dma_status[63:56];
assign builder_genericstandalone_csrbank7_dma_byte_count6_w = main_rtio_analyzer_dma_status[55:48];
assign builder_genericstandalone_csrbank7_dma_byte_count5_w = main_rtio_analyzer_dma_status[47:40];
assign builder_genericstandalone_csrbank7_dma_byte_count4_w = main_rtio_analyzer_dma_status[39:32];
assign builder_genericstandalone_csrbank7_dma_byte_count3_w = main_rtio_analyzer_dma_status[31:24];
assign builder_genericstandalone_csrbank7_dma_byte_count2_w = main_rtio_analyzer_dma_status[23:16];
assign builder_genericstandalone_csrbank7_dma_byte_count1_w = main_rtio_analyzer_dma_status[15:8];
assign builder_genericstandalone_csrbank7_dma_byte_count0_w = main_rtio_analyzer_dma_status[7:0];
assign builder_genericstandalone_csrbank8_sel = (builder_genericstandalone_interface8_bank_bus_adr[13:9] == 4'd15);
assign main_rtio_core_reset_r = builder_genericstandalone_interface8_bank_bus_dat_w[0];
assign main_rtio_core_reset_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 1'd0));
assign main_rtio_core_reset_phy_r = builder_genericstandalone_interface8_bank_bus_dat_w[0];
assign main_rtio_core_reset_phy_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 1'd1));
assign main_rtio_core_async_error_r = builder_genericstandalone_interface8_bank_bus_dat_w[2:0];
assign main_rtio_core_async_error_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 2'd2));
assign builder_genericstandalone_csrbank8_collision_channel1_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_collision_channel1_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 2'd3));
assign builder_genericstandalone_csrbank8_collision_channel0_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_collision_channel0_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 3'd4));
assign builder_genericstandalone_csrbank8_busy_channel1_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_busy_channel1_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 3'd5));
assign builder_genericstandalone_csrbank8_busy_channel0_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_busy_channel0_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 3'd6));
assign builder_genericstandalone_csrbank8_sequence_error_channel1_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_sequence_error_channel1_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 3'd7));
assign builder_genericstandalone_csrbank8_sequence_error_channel0_r = builder_genericstandalone_interface8_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank8_sequence_error_channel0_re = ((builder_genericstandalone_csrbank8_sel & builder_genericstandalone_interface8_bank_bus_we) & (builder_genericstandalone_interface8_bank_bus_adr[3:0] == 4'd8));
assign builder_genericstandalone_csrbank8_collision_channel1_w = main_rtio_core_collision_channel_status[15:8];
assign builder_genericstandalone_csrbank8_collision_channel0_w = main_rtio_core_collision_channel_status[7:0];
assign builder_genericstandalone_csrbank8_busy_channel1_w = main_rtio_core_busy_channel_status[15:8];
assign builder_genericstandalone_csrbank8_busy_channel0_w = main_rtio_core_busy_channel_status[7:0];
assign builder_genericstandalone_csrbank8_sequence_error_channel1_w = main_rtio_core_sequence_error_channel_status[15:8];
assign builder_genericstandalone_csrbank8_sequence_error_channel0_w = main_rtio_core_sequence_error_channel_status[7:0];
assign builder_genericstandalone_csrbank9_sel = (builder_genericstandalone_interface9_bank_bus_adr[13:9] == 4'd14);
assign builder_genericstandalone_csrbank9_pll_reset0_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_pll_reset0_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[0] == 1'd0));
assign builder_genericstandalone_csrbank9_pll_locked_r = builder_genericstandalone_interface9_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank9_pll_locked_re = ((builder_genericstandalone_csrbank9_sel & builder_genericstandalone_interface9_bank_bus_we) & (builder_genericstandalone_interface9_bank_bus_adr[0] == 1'd1));
assign main_rtio_crg_storage = main_rtio_crg_storage_full;
assign builder_genericstandalone_csrbank9_pll_reset0_w = main_rtio_crg_storage_full;
assign builder_genericstandalone_csrbank9_pll_locked_w = main_rtio_crg_pll_locked_status;
assign builder_genericstandalone_csrbank10_sel = (builder_genericstandalone_interface10_bank_bus_adr[13:9] == 5'd16);
assign builder_genericstandalone_csrbank10_mon_chan_sel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank10_mon_chan_sel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 1'd0));
assign builder_genericstandalone_csrbank10_mon_probe_sel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank10_mon_probe_sel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 1'd1));
assign main_mon_value_update_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign main_mon_value_update_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 2'd2));
assign builder_genericstandalone_csrbank10_mon_value_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank10_mon_value_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 2'd3));
assign builder_genericstandalone_csrbank10_inj_chan_sel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank10_inj_chan_sel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 3'd4));
assign builder_genericstandalone_csrbank10_inj_override_sel0_r = builder_genericstandalone_interface10_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank10_inj_override_sel0_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 3'd5));
assign main_inj_value_r = builder_genericstandalone_interface10_bank_bus_dat_w[0];
assign main_inj_value_re = ((builder_genericstandalone_csrbank10_sel & builder_genericstandalone_interface10_bank_bus_we) & (builder_genericstandalone_interface10_bank_bus_adr[2:0] == 3'd6));
assign main_mon_chan_sel_storage = main_mon_chan_sel_storage_full[5:0];
assign builder_genericstandalone_csrbank10_mon_chan_sel0_w = main_mon_chan_sel_storage_full[5:0];
assign main_mon_probe_sel_storage = main_mon_probe_sel_storage_full;
assign builder_genericstandalone_csrbank10_mon_probe_sel0_w = main_mon_probe_sel_storage_full;
assign builder_genericstandalone_csrbank10_mon_value_w = main_mon_status;
assign main_inj_chan_sel_storage = main_inj_chan_sel_storage_full[5:0];
assign builder_genericstandalone_csrbank10_inj_chan_sel0_w = main_inj_chan_sel_storage_full[5:0];
assign main_inj_override_sel_storage = main_inj_override_sel_storage_full[1:0];
assign builder_genericstandalone_csrbank10_inj_override_sel0_w = main_inj_override_sel_storage_full[1:0];
assign builder_genericstandalone_csrbank11_sel = (builder_genericstandalone_interface11_bank_bus_adr[13:9] == 4'd8);
assign builder_genericstandalone_csrbank11_bitbang0_r = builder_genericstandalone_interface11_bank_bus_dat_w[3:0];
assign builder_genericstandalone_csrbank11_bitbang0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank11_miso_r = builder_genericstandalone_interface11_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank11_miso_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank11_bitbang_en0_r = builder_genericstandalone_interface11_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank11_bitbang_en0_re = ((builder_genericstandalone_csrbank11_sel & builder_genericstandalone_interface11_bank_bus_we) & (builder_genericstandalone_interface11_bank_bus_adr[1:0] == 2'd2));
assign main_genericstandalone_genericstandalone_spiflash_bitbang_storage = main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0];
assign builder_genericstandalone_csrbank11_bitbang0_w = main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0];
assign builder_genericstandalone_csrbank11_miso_w = main_genericstandalone_genericstandalone_spiflash_status;
assign main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage = main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full;
assign builder_genericstandalone_csrbank11_bitbang_en0_w = main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full;
assign builder_genericstandalone_csrbank12_sel = (builder_genericstandalone_interface12_bank_bus_adr[13:9] == 2'd3);
assign builder_genericstandalone_csrbank12_load7_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load7_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 1'd0));
assign builder_genericstandalone_csrbank12_load6_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load6_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 1'd1));
assign builder_genericstandalone_csrbank12_load5_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load5_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 2'd2));
assign builder_genericstandalone_csrbank12_load4_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load4_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 2'd3));
assign builder_genericstandalone_csrbank12_load3_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load3_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 3'd4));
assign builder_genericstandalone_csrbank12_load2_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load2_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 3'd5));
assign builder_genericstandalone_csrbank12_load1_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load1_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 3'd6));
assign builder_genericstandalone_csrbank12_load0_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_load0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 3'd7));
assign builder_genericstandalone_csrbank12_reload7_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload7_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd8));
assign builder_genericstandalone_csrbank12_reload6_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload6_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd9));
assign builder_genericstandalone_csrbank12_reload5_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload5_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd10));
assign builder_genericstandalone_csrbank12_reload4_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload4_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd11));
assign builder_genericstandalone_csrbank12_reload3_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload3_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd12));
assign builder_genericstandalone_csrbank12_reload2_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload2_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd13));
assign builder_genericstandalone_csrbank12_reload1_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload1_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd14));
assign builder_genericstandalone_csrbank12_reload0_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_reload0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 4'd15));
assign builder_genericstandalone_csrbank12_en0_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank12_en0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd16));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd17));
assign builder_genericstandalone_csrbank12_value7_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value7_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd18));
assign builder_genericstandalone_csrbank12_value6_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value6_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd19));
assign builder_genericstandalone_csrbank12_value5_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value5_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd20));
assign builder_genericstandalone_csrbank12_value4_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value4_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd21));
assign builder_genericstandalone_csrbank12_value3_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value3_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd22));
assign builder_genericstandalone_csrbank12_value2_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value2_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd23));
assign builder_genericstandalone_csrbank12_value1_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value1_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd24));
assign builder_genericstandalone_csrbank12_value0_r = builder_genericstandalone_interface12_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank12_value0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd25));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd26));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd27));
assign builder_genericstandalone_csrbank12_ev_enable0_r = builder_genericstandalone_interface12_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank12_ev_enable0_re = ((builder_genericstandalone_csrbank12_sel & builder_genericstandalone_interface12_bank_bus_we) & (builder_genericstandalone_interface12_bank_bus_adr[4:0] == 5'd28));
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:0];
assign builder_genericstandalone_csrbank12_load7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:56];
assign builder_genericstandalone_csrbank12_load6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[55:48];
assign builder_genericstandalone_csrbank12_load5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[47:40];
assign builder_genericstandalone_csrbank12_load4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[39:32];
assign builder_genericstandalone_csrbank12_load3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[31:24];
assign builder_genericstandalone_csrbank12_load2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[23:16];
assign builder_genericstandalone_csrbank12_load1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[15:8];
assign builder_genericstandalone_csrbank12_load0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:0];
assign builder_genericstandalone_csrbank12_reload7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:56];
assign builder_genericstandalone_csrbank12_reload6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[55:48];
assign builder_genericstandalone_csrbank12_reload5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[47:40];
assign builder_genericstandalone_csrbank12_reload4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[39:32];
assign builder_genericstandalone_csrbank12_reload3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[31:24];
assign builder_genericstandalone_csrbank12_reload2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[23:16];
assign builder_genericstandalone_csrbank12_reload1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[15:8];
assign builder_genericstandalone_csrbank12_reload0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full;
assign builder_genericstandalone_csrbank12_en0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full;
assign builder_genericstandalone_csrbank12_value7_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[63:56];
assign builder_genericstandalone_csrbank12_value6_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[55:48];
assign builder_genericstandalone_csrbank12_value5_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[47:40];
assign builder_genericstandalone_csrbank12_value4_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[39:32];
assign builder_genericstandalone_csrbank12_value3_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[31:24];
assign builder_genericstandalone_csrbank12_value2_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[23:16];
assign builder_genericstandalone_csrbank12_value1_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[15:8];
assign builder_genericstandalone_csrbank12_value0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage = main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full;
assign builder_genericstandalone_csrbank12_ev_enable0_w = main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full;
assign builder_genericstandalone_csrbank13_sel = (builder_genericstandalone_interface13_bank_bus_adr[13:9] == 3'd4);
assign builder_genericstandalone_csrbank13_enable_null0_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank13_enable_null0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 1'd0));
assign builder_genericstandalone_csrbank13_enable_prog0_r = builder_genericstandalone_interface13_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank13_enable_prog0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 1'd1));
assign builder_genericstandalone_csrbank13_prog_address3_r = builder_genericstandalone_interface13_bank_bus_dat_w[5:0];
assign builder_genericstandalone_csrbank13_prog_address3_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 2'd2));
assign builder_genericstandalone_csrbank13_prog_address2_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_prog_address2_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 2'd3));
assign builder_genericstandalone_csrbank13_prog_address1_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_prog_address1_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 3'd4));
assign builder_genericstandalone_csrbank13_prog_address0_r = builder_genericstandalone_interface13_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank13_prog_address0_re = ((builder_genericstandalone_csrbank13_sel & builder_genericstandalone_interface13_bank_bus_we) & (builder_genericstandalone_interface13_bank_bus_adr[2:0] == 3'd5));
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage = main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage_full;
assign builder_genericstandalone_csrbank13_enable_null0_w = main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage_full;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage = main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage_full;
assign builder_genericstandalone_csrbank13_enable_prog0_w = main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage_full;
assign main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage = main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[29:12];
assign builder_genericstandalone_csrbank13_prog_address3_w = main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[29:24];
assign builder_genericstandalone_csrbank13_prog_address2_w = main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[23:16];
assign builder_genericstandalone_csrbank13_prog_address1_w = {main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[15:12], {4{1'd0}}};
assign builder_genericstandalone_csrbank13_prog_address0_w = 1'd0;
assign builder_genericstandalone_csrbank14_sel = (builder_genericstandalone_interface14_bank_bus_adr[13:9] == 1'd1);
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_r = builder_genericstandalone_interface14_bank_bus_dat_w[7:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 1'd0));
assign builder_genericstandalone_csrbank14_txfull_r = builder_genericstandalone_interface14_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank14_txfull_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 1'd1));
assign builder_genericstandalone_csrbank14_rxempty_r = builder_genericstandalone_interface14_bank_bus_dat_w[0];
assign builder_genericstandalone_csrbank14_rxempty_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 2'd2));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_status_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_status_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 2'd3));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_pending_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign main_genericstandalone_genericstandalone_genericstandalone_uart_pending_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 3'd4));
assign builder_genericstandalone_csrbank14_ev_enable0_r = builder_genericstandalone_interface14_bank_bus_dat_w[1:0];
assign builder_genericstandalone_csrbank14_ev_enable0_re = ((builder_genericstandalone_csrbank14_sel & builder_genericstandalone_interface14_bank_bus_we) & (builder_genericstandalone_interface14_bank_bus_adr[2:0] == 3'd5));
assign builder_genericstandalone_csrbank14_txfull_w = main_genericstandalone_genericstandalone_genericstandalone_uart_txfull_status;
assign builder_genericstandalone_csrbank14_rxempty_w = main_genericstandalone_genericstandalone_genericstandalone_uart_rxempty_status;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_storage = main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0];
assign builder_genericstandalone_csrbank14_ev_enable0_w = main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0];
assign builder_genericstandalone_csrbank15_sel = (builder_genericstandalone_interface15_bank_bus_adr[13:9] == 1'd0);
assign builder_genericstandalone_csrbank15_tuning_word3_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word3_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 1'd0));
assign builder_genericstandalone_csrbank15_tuning_word2_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word2_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 1'd1));
assign builder_genericstandalone_csrbank15_tuning_word1_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word1_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 2'd2));
assign builder_genericstandalone_csrbank15_tuning_word0_r = builder_genericstandalone_interface15_bank_bus_dat_w[7:0];
assign builder_genericstandalone_csrbank15_tuning_word0_re = ((builder_genericstandalone_csrbank15_sel & builder_genericstandalone_interface15_bank_bus_we) & (builder_genericstandalone_interface15_bank_bus_adr[1:0] == 2'd3));
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:0];
assign builder_genericstandalone_csrbank15_tuning_word3_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:24];
assign builder_genericstandalone_csrbank15_tuning_word2_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[23:16];
assign builder_genericstandalone_csrbank15_tuning_word1_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[15:8];
assign builder_genericstandalone_csrbank15_tuning_word0_w = main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[7:0];
assign builder_genericstandalone_interface0_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface1_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface2_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface3_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface4_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface5_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface6_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface7_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface8_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface9_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface10_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface11_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface12_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface13_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface14_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface15_bank_bus_adr = main_genericstandalone_genericstandalone_genericstandalone_interface_adr;
assign builder_genericstandalone_interface0_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface1_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface2_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface3_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface4_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface5_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface6_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface7_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface8_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface9_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface10_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface11_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface12_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface13_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface14_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface15_bank_bus_we = main_genericstandalone_genericstandalone_genericstandalone_interface_we;
assign builder_genericstandalone_interface0_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface1_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface2_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface3_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface4_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface5_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface6_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface7_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface8_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface9_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface10_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface11_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface12_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface13_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface14_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign builder_genericstandalone_interface15_bank_bus_dat_w = main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w;
assign main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r = (((((((((((((((builder_genericstandalone_interface0_bank_bus_dat_r | builder_genericstandalone_interface1_bank_bus_dat_r) | builder_genericstandalone_interface2_bank_bus_dat_r) | builder_genericstandalone_interface3_bank_bus_dat_r) | builder_genericstandalone_interface4_bank_bus_dat_r) | builder_genericstandalone_interface5_bank_bus_dat_r) | builder_genericstandalone_interface6_bank_bus_dat_r) | builder_genericstandalone_interface7_bank_bus_dat_r) | builder_genericstandalone_interface8_bank_bus_dat_r) | builder_genericstandalone_interface9_bank_bus_dat_r) | builder_genericstandalone_interface10_bank_bus_dat_r) | builder_genericstandalone_interface11_bank_bus_dat_r) | builder_genericstandalone_interface12_bank_bus_dat_r) | builder_genericstandalone_interface13_bank_bus_dat_r) | builder_genericstandalone_interface14_bank_bus_dat_r) | builder_genericstandalone_interface15_bank_bus_dat_r);

// synthesis translate_off
reg dummy_d_168;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed0 <= 30'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed0 <= main_genericstandalone_kernel_cpu_ibus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed0 <= main_genericstandalone_kernel_cpu_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_168 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_169;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed1 <= 32'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed1 <= main_genericstandalone_kernel_cpu_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed1 <= main_genericstandalone_kernel_cpu_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_169 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_170;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed2 <= 4'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed2 <= main_genericstandalone_kernel_cpu_ibus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed2 <= main_genericstandalone_kernel_cpu_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_170 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_171;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed3 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed3 <= main_genericstandalone_kernel_cpu_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed3 <= main_genericstandalone_kernel_cpu_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_171 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_172;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed4 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed4 <= main_genericstandalone_kernel_cpu_ibus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed4 <= main_genericstandalone_kernel_cpu_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_172 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_173;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed5 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed5 <= main_genericstandalone_kernel_cpu_ibus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed5 <= main_genericstandalone_kernel_cpu_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_173 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_174;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed6 <= 3'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed6 <= main_genericstandalone_kernel_cpu_ibus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed6 <= main_genericstandalone_kernel_cpu_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_174 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_175;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed7 <= 2'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed7 <= main_genericstandalone_kernel_cpu_ibus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed7 <= main_genericstandalone_kernel_cpu_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_175 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_176;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed8 <= 1'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record0_writable;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record1_writable;
		end
		2'd2: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record2_writable;
		end
		2'd3: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record3_writable;
		end
		3'd4: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record4_writable;
		end
		3'd5: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record5_writable;
		end
		3'd6: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record6_writable;
		end
		default: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record7_writable;
		end
	endcase
// synthesis translate_off
	dummy_d_176 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_177;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed9 <= 2'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow0, (main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & (~main_rtio_core_inputs_overflow0))};
		end
		1'd1: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow1, (main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & (~main_rtio_core_inputs_overflow1))};
		end
		2'd2: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow2, (main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & (~main_rtio_core_inputs_overflow2))};
		end
		2'd3: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow3, (main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & (~main_rtio_core_inputs_overflow3))};
		end
		3'd4: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow4, (main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & (~main_rtio_core_inputs_overflow4))};
		end
		3'd5: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow5, (main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & (~main_rtio_core_inputs_overflow5))};
		end
		3'd6: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow6, (main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & (~main_rtio_core_inputs_overflow6))};
		end
		3'd7: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow7, (main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable & (~main_rtio_core_inputs_overflow7))};
		end
		4'd8: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd9: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd10: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd11: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd12: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd13: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd14: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd15: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd16: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow8, (main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable & (~main_rtio_core_inputs_overflow8))};
		end
		5'd17: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd18: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd19: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd20: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd21: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd22: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow9, (main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable & (~main_rtio_core_inputs_overflow9))};
		end
		5'd23: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd24: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd25: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd26: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd27: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd28: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow10, (main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable & (~main_rtio_core_inputs_overflow10))};
		end
		5'd29: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd30: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd31: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd32: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd33: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd34: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd35: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_177 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_178;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed10 <= 2'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed10 <= main_rtio_cri_cmd;
		end
		default: begin
			builder_comb_rhs_array_muxed10 <= main_dma_cri_master_cri_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_178 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_179;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed11 <= 24'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed11 <= main_rtio_cri_chan_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed11 <= main_dma_cri_master_cri_chan_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_179 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_180;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed12 <= 64'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed12 <= main_rtio_cri_o_timestamp;
		end
		default: begin
			builder_comb_rhs_array_muxed12 <= main_dma_cri_master_cri_o_timestamp;
		end
	endcase
// synthesis translate_off
	dummy_d_180 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_181;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed13 <= 512'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed13 <= main_rtio_cri_o_data;
		end
		default: begin
			builder_comb_rhs_array_muxed13 <= main_dma_cri_master_cri_o_data;
		end
	endcase
// synthesis translate_off
	dummy_d_181 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_182;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed14 <= 8'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed14 <= main_rtio_cri_o_address;
		end
		default: begin
			builder_comb_rhs_array_muxed14 <= main_dma_cri_master_cri_o_address;
		end
	endcase
// synthesis translate_off
	dummy_d_182 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_183;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed15 <= 64'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed15 <= main_rtio_cri_i_timeout;
		end
		default: begin
			builder_comb_rhs_array_muxed15 <= main_dma_cri_master_cri_i_timeout;
		end
	endcase
// synthesis translate_off
	dummy_d_183 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_184;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed17 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed17 <= main_inj_o_sys0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed17 <= main_inj_o_sys1;
		end
		default: begin
			builder_comb_rhs_array_muxed17 <= main_inj_o_sys2;
		end
	endcase
// synthesis translate_off
	dummy_d_184 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_185;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed18 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed18 <= main_inj_o_sys3;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed18 <= main_inj_o_sys4;
		end
		default: begin
			builder_comb_rhs_array_muxed18 <= main_inj_o_sys5;
		end
	endcase
// synthesis translate_off
	dummy_d_185 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_186;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed19 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed19 <= main_inj_o_sys6;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed19 <= main_inj_o_sys7;
		end
		default: begin
			builder_comb_rhs_array_muxed19 <= main_inj_o_sys8;
		end
	endcase
// synthesis translate_off
	dummy_d_186 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_187;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed20 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys9;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys10;
		end
		default: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys11;
		end
	endcase
// synthesis translate_off
	dummy_d_187 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_188;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed21 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed21 <= main_inj_o_sys12;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed21 <= main_inj_o_sys13;
		end
		default: begin
			builder_comb_rhs_array_muxed21 <= main_inj_o_sys14;
		end
	endcase
// synthesis translate_off
	dummy_d_188 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_189;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed22 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed22 <= main_inj_o_sys15;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed22 <= main_inj_o_sys16;
		end
		default: begin
			builder_comb_rhs_array_muxed22 <= main_inj_o_sys17;
		end
	endcase
// synthesis translate_off
	dummy_d_189 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_190;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed23 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed23 <= main_inj_o_sys18;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed23 <= main_inj_o_sys19;
		end
		default: begin
			builder_comb_rhs_array_muxed23 <= main_inj_o_sys20;
		end
	endcase
// synthesis translate_off
	dummy_d_190 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_191;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed24 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys21;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys22;
		end
		default: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys23;
		end
	endcase
// synthesis translate_off
	dummy_d_191 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_192;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed25 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed25 <= main_inj_o_sys24;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed25 <= main_inj_o_sys25;
		end
		default: begin
			builder_comb_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_192 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_193;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed26 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed26 <= main_inj_o_sys26;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed26 <= main_inj_o_sys27;
		end
		default: begin
			builder_comb_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_193 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_194;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed27 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed27 <= main_inj_o_sys28;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed27 <= main_inj_o_sys29;
		end
		default: begin
			builder_comb_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_194 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_195;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed28 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed28 <= main_inj_o_sys30;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed28 <= main_inj_o_sys31;
		end
		default: begin
			builder_comb_rhs_array_muxed28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_195 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_196;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed29 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed29 <= main_inj_o_sys32;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed29 <= main_inj_o_sys33;
		end
		default: begin
			builder_comb_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_196 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_197;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed30 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed30 <= main_inj_o_sys34;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed30 <= main_inj_o_sys35;
		end
		default: begin
			builder_comb_rhs_array_muxed30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_197 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_198;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed31 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed31 <= main_inj_o_sys36;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed31 <= main_inj_o_sys37;
		end
		default: begin
			builder_comb_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_198 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_199;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed32 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed32 <= main_inj_o_sys38;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed32 <= main_inj_o_sys39;
		end
		default: begin
			builder_comb_rhs_array_muxed32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_199 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_200;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed33 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed33 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed33 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_200 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_201;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed34 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed34 <= main_inj_o_sys40;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed34 <= main_inj_o_sys41;
		end
		default: begin
			builder_comb_rhs_array_muxed34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_201 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_202;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed35 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed35 <= main_inj_o_sys42;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed35 <= main_inj_o_sys43;
		end
		default: begin
			builder_comb_rhs_array_muxed35 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_202 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_203;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed36 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed36 <= main_inj_o_sys44;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed36 <= main_inj_o_sys45;
		end
		default: begin
			builder_comb_rhs_array_muxed36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_203 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_204;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed37 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed37 <= main_inj_o_sys46;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed37 <= main_inj_o_sys47;
		end
		default: begin
			builder_comb_rhs_array_muxed37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_204 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_205;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed38 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed38 <= main_inj_o_sys48;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed38 <= main_inj_o_sys49;
		end
		default: begin
			builder_comb_rhs_array_muxed38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_205 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_206;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed39 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_206 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_207;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed40 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed40 <= main_inj_o_sys50;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed40 <= main_inj_o_sys51;
		end
		default: begin
			builder_comb_rhs_array_muxed40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_207 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_208;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed41 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed41 <= main_inj_o_sys52;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed41 <= main_inj_o_sys53;
		end
		default: begin
			builder_comb_rhs_array_muxed41 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_208 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_209;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed42 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed42 <= main_inj_o_sys54;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed42 <= main_inj_o_sys55;
		end
		default: begin
			builder_comb_rhs_array_muxed42 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_209 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_210;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed43 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed43 <= main_inj_o_sys56;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed43 <= main_inj_o_sys57;
		end
		default: begin
			builder_comb_rhs_array_muxed43 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_210 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_211;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed44 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed44 <= main_inj_o_sys58;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed44 <= main_inj_o_sys59;
		end
		default: begin
			builder_comb_rhs_array_muxed44 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_211 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_212;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed45 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_212 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_213;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed46 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed46 <= main_inj_o_sys60;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed46 <= main_inj_o_sys61;
		end
		default: begin
			builder_comb_rhs_array_muxed46 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_213 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_214;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed47 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed47 <= main_inj_o_sys62;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed47 <= main_inj_o_sys63;
		end
		default: begin
			builder_comb_rhs_array_muxed47 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_214 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_215;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed48 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed48 <= main_inj_o_sys64;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed48 <= main_inj_o_sys65;
		end
		default: begin
			builder_comb_rhs_array_muxed48 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_215 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_216;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed49 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed49 <= main_inj_o_sys66;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed49 <= main_inj_o_sys67;
		end
		default: begin
			builder_comb_rhs_array_muxed49 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_216 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_217;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed50 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed50 <= main_inj_o_sys68;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed50 <= main_inj_o_sys69;
		end
		default: begin
			builder_comb_rhs_array_muxed50 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_217 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_218;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed51 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed51 <= main_inj_o_sys70;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed51 <= main_inj_o_sys71;
		end
		default: begin
			builder_comb_rhs_array_muxed51 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_218 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_219;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed52 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed52 <= main_inj_o_sys72;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed52 <= main_inj_o_sys73;
		end
		default: begin
			builder_comb_rhs_array_muxed52 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_219 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_220;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed53 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed53 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed53 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed53 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_220 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_221;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed16 <= 1'd0;
	case (main_inj_chan_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed17;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed18;
		end
		2'd2: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed19;
		end
		2'd3: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed20;
		end
		3'd4: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed21;
		end
		3'd5: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed22;
		end
		3'd6: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed23;
		end
		3'd7: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed24;
		end
		4'd8: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed25;
		end
		4'd9: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed26;
		end
		4'd10: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed27;
		end
		4'd11: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed28;
		end
		4'd12: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed29;
		end
		4'd13: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed30;
		end
		4'd14: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed31;
		end
		4'd15: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed32;
		end
		5'd16: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed33;
		end
		5'd17: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed34;
		end
		5'd18: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed35;
		end
		5'd19: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed36;
		end
		5'd20: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed37;
		end
		5'd21: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed38;
		end
		5'd22: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed39;
		end
		5'd23: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed40;
		end
		5'd24: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed41;
		end
		5'd25: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed42;
		end
		5'd26: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed43;
		end
		5'd27: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed44;
		end
		5'd28: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed45;
		end
		5'd29: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed46;
		end
		5'd30: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed47;
		end
		5'd31: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed48;
		end
		6'd32: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed49;
		end
		6'd33: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed50;
		end
		6'd34: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed51;
		end
		6'd35: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed52;
		end
		default: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed53;
		end
	endcase
// synthesis translate_off
	dummy_d_221 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_222;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed54 <= 30'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed54 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed54 <= main_genericstandalone_kernel_cpu_wb_sdram_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_222 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_223;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed55 <= 32'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed55 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed55 <= main_genericstandalone_kernel_cpu_wb_sdram_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_223 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_224;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed56 <= 4'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed56 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed56 <= main_genericstandalone_kernel_cpu_wb_sdram_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_224 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_225;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed57 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed57 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed57 <= main_genericstandalone_kernel_cpu_wb_sdram_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_225 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_226;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed58 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed58 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed58 <= main_genericstandalone_kernel_cpu_wb_sdram_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_226 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_227;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed59 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed59 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_we;
		end
		default: begin
			builder_comb_rhs_array_muxed59 <= main_genericstandalone_kernel_cpu_wb_sdram_we;
		end
	endcase
// synthesis translate_off
	dummy_d_227 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_228;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed60 <= 3'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed60 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed60 <= main_genericstandalone_kernel_cpu_wb_sdram_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_228 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_229;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed61 <= 2'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed61 <= main_genericstandalone_genericstandalone_genericstandalone_wb_sdram_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed61 <= main_genericstandalone_kernel_cpu_wb_sdram_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_229 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_230;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed62 <= 30'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed62 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_adr;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed62 <= main_genericstandalone_interface0_bus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed62 <= main_genericstandalone_interface1_bus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_230 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_231;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed63 <= 128'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed63 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_dat_w;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed63 <= main_genericstandalone_interface0_bus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed63 <= main_genericstandalone_interface1_bus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_231 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_232;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed64 <= 16'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed64 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_sel;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed64 <= main_genericstandalone_interface0_bus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed64 <= main_genericstandalone_interface1_bus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_232 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_233;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed65 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed65 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cyc;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed65 <= main_genericstandalone_interface0_bus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed65 <= main_genericstandalone_interface1_bus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_233 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_234;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed66 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed66 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_stb;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed66 <= main_genericstandalone_interface0_bus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed66 <= main_genericstandalone_interface1_bus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_234 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_235;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed67 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed67 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_we;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed67 <= main_genericstandalone_interface0_bus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed67 <= main_genericstandalone_interface1_bus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_235 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_236;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed68 <= 3'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed68 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_cti;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed68 <= main_genericstandalone_interface0_bus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed68 <= main_genericstandalone_interface1_bus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_236 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_237;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed69 <= 2'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed69 <= main_genericstandalone_genericstandalone_genericstandalone_bridge_if_bus_bte;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed69 <= main_genericstandalone_interface0_bus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed69 <= main_genericstandalone_interface1_bus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_237 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_238;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed70 <= 30'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed70 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed70 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_238 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_239;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed71 <= 32'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed71 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed71 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_239 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_240;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed72 <= 4'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed72 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed72 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_240 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_241;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed73 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed73 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed73 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_241 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_242;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed74 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed74 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed74 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_242 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_243;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed75 <= 1'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed75 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed75 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_we;
		end
	endcase
// synthesis translate_off
	dummy_d_243 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_244;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed76 <= 3'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed76 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed76 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_244 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_245;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed77 <= 2'd0;
	case (builder_genericstandalone_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed77 <= main_genericstandalone_genericstandalone_genericstandalone_ibus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed77 <= main_genericstandalone_genericstandalone_genericstandalone_tmpu_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_245 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_246;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed0 <= 3'd4;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed0 <= 2'd3;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed0 <= 2'd2;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed0 <= 3'd6;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed0 <= 3'd7;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd1;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed0 <= 3'd5;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_246 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_247;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed0 <= 3'd5;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed0 <= 1'd1;
		end
		3'd7: begin
			builder_sync_f_t_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		4'd9: begin
			builder_sync_f_t_array_muxed0 <= 3'd6;
		end
		4'd10: begin
			builder_sync_f_t_array_muxed0 <= 2'd2;
		end
		4'd11: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_t_array_muxed0 <= 2'd3;
		end
		4'd13: begin
			builder_sync_f_t_array_muxed0 <= 3'd4;
		end
		4'd14: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
		default: begin
			builder_sync_f_t_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_247 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_248;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_array_muxed0 <= 3'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			builder_sync_f_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd7;
		end
		2'd2: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd4;
		end
		2'd3: begin
			builder_sync_f_rhs_array_muxed0 <= 2'd3;
		end
		3'd4: begin
			builder_sync_f_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_f_rhs_array_muxed0 <= 2'd2;
		end
		3'd6: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd6;
		end
		3'd7: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd7;
		end
		4'd9: begin
			builder_sync_f_rhs_array_muxed0 <= 1'd1;
		end
		4'd10: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd5;
		end
		4'd11: begin
			builder_sync_f_rhs_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_array_muxed0 <= 2'd3;
		end
		4'd13: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd4;
		end
		4'd14: begin
			builder_sync_f_rhs_array_muxed0 <= 3'd7;
		end
		default: begin
			builder_sync_f_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_248 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_249;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed0 <= 5'd0;
	case (main_genericstandalone_pcs_receivepath_input_msb_first[9:4])
		1'd0: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed0 <= 5'd23;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed0 <= 4'd8;
		end
		3'd7: begin
			builder_sync_rhs_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		4'd9: begin
			builder_sync_rhs_array_muxed0 <= 5'd27;
		end
		4'd10: begin
			builder_sync_rhs_array_muxed0 <= 3'd4;
		end
		4'd11: begin
			builder_sync_rhs_array_muxed0 <= 5'd20;
		end
		4'd12: begin
			builder_sync_rhs_array_muxed0 <= 5'd24;
		end
		4'd13: begin
			builder_sync_rhs_array_muxed0 <= 4'd12;
		end
		4'd14: begin
			builder_sync_rhs_array_muxed0 <= 5'd28;
		end
		4'd15: begin
			builder_sync_rhs_array_muxed0 <= 5'd28;
		end
		5'd16: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		5'd17: begin
			builder_sync_rhs_array_muxed0 <= 5'd29;
		end
		5'd18: begin
			builder_sync_rhs_array_muxed0 <= 2'd2;
		end
		5'd19: begin
			builder_sync_rhs_array_muxed0 <= 5'd18;
		end
		5'd20: begin
			builder_sync_rhs_array_muxed0 <= 5'd31;
		end
		5'd21: begin
			builder_sync_rhs_array_muxed0 <= 4'd10;
		end
		5'd22: begin
			builder_sync_rhs_array_muxed0 <= 5'd26;
		end
		5'd23: begin
			builder_sync_rhs_array_muxed0 <= 4'd15;
		end
		5'd24: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		5'd25: begin
			builder_sync_rhs_array_muxed0 <= 3'd6;
		end
		5'd26: begin
			builder_sync_rhs_array_muxed0 <= 5'd22;
		end
		5'd27: begin
			builder_sync_rhs_array_muxed0 <= 5'd16;
		end
		5'd28: begin
			builder_sync_rhs_array_muxed0 <= 4'd14;
		end
		5'd29: begin
			builder_sync_rhs_array_muxed0 <= 1'd1;
		end
		5'd30: begin
			builder_sync_rhs_array_muxed0 <= 5'd30;
		end
		5'd31: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd32: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd33: begin
			builder_sync_rhs_array_muxed0 <= 5'd30;
		end
		6'd34: begin
			builder_sync_rhs_array_muxed0 <= 1'd1;
		end
		6'd35: begin
			builder_sync_rhs_array_muxed0 <= 5'd17;
		end
		6'd36: begin
			builder_sync_rhs_array_muxed0 <= 5'd16;
		end
		6'd37: begin
			builder_sync_rhs_array_muxed0 <= 4'd9;
		end
		6'd38: begin
			builder_sync_rhs_array_muxed0 <= 5'd25;
		end
		6'd39: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd40: begin
			builder_sync_rhs_array_muxed0 <= 4'd15;
		end
		6'd41: begin
			builder_sync_rhs_array_muxed0 <= 3'd5;
		end
		6'd42: begin
			builder_sync_rhs_array_muxed0 <= 5'd21;
		end
		6'd43: begin
			builder_sync_rhs_array_muxed0 <= 5'd31;
		end
		6'd44: begin
			builder_sync_rhs_array_muxed0 <= 4'd13;
		end
		6'd45: begin
			builder_sync_rhs_array_muxed0 <= 2'd2;
		end
		6'd46: begin
			builder_sync_rhs_array_muxed0 <= 5'd29;
		end
		6'd47: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd48: begin
			builder_sync_rhs_array_muxed0 <= 5'd28;
		end
		6'd49: begin
			builder_sync_rhs_array_muxed0 <= 2'd3;
		end
		6'd50: begin
			builder_sync_rhs_array_muxed0 <= 5'd19;
		end
		6'd51: begin
			builder_sync_rhs_array_muxed0 <= 5'd24;
		end
		6'd52: begin
			builder_sync_rhs_array_muxed0 <= 4'd11;
		end
		6'd53: begin
			builder_sync_rhs_array_muxed0 <= 3'd4;
		end
		6'd54: begin
			builder_sync_rhs_array_muxed0 <= 5'd27;
		end
		6'd55: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd56: begin
			builder_sync_rhs_array_muxed0 <= 3'd7;
		end
		6'd57: begin
			builder_sync_rhs_array_muxed0 <= 4'd8;
		end
		6'd58: begin
			builder_sync_rhs_array_muxed0 <= 5'd23;
		end
		6'd59: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd60: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd61: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd62: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
		default: begin
			builder_sync_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_249 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_250;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_array_muxed1 <= 6'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[4:0])
		1'd0: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd24;
		end
		1'd1: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd34;
		end
		2'd2: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd18;
		end
		2'd3: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd49;
		end
		3'd4: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd10;
		end
		3'd5: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd41;
		end
		3'd6: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd25;
		end
		3'd7: begin
			builder_sync_f_rhs_array_muxed1 <= 3'd7;
		end
		4'd8: begin
			builder_sync_f_rhs_array_muxed1 <= 3'd6;
		end
		4'd9: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd37;
		end
		4'd10: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd21;
		end
		4'd11: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd52;
		end
		4'd12: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd13;
		end
		4'd13: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd44;
		end
		4'd14: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd28;
		end
		4'd15: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd40;
		end
		5'd16: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd36;
		end
		5'd17: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd35;
		end
		5'd18: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd19;
		end
		5'd19: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd50;
		end
		5'd20: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd11;
		end
		5'd21: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd42;
		end
		5'd22: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd26;
		end
		5'd23: begin
			builder_sync_f_rhs_array_muxed1 <= 3'd5;
		end
		5'd24: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd12;
		end
		5'd25: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd38;
		end
		5'd26: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd22;
		end
		5'd27: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd9;
		end
		5'd28: begin
			builder_sync_f_rhs_array_muxed1 <= 4'd14;
		end
		5'd29: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd17;
		end
		5'd30: begin
			builder_sync_f_rhs_array_muxed1 <= 6'd33;
		end
		default: begin
			builder_sync_f_rhs_array_muxed1 <= 5'd20;
		end
	endcase
// synthesis translate_off
	dummy_d_250 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_251;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_array_muxed2 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[4:0])
		1'd0: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		2'd3: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd7: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd8: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		4'd9: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd10: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd11: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd13: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd14: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd15: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd16: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd17: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd18: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd19: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd20: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd21: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd22: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd23: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd24: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd25: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd26: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd27: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd28: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd29: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd30: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
		default: begin
			builder_sync_f_rhs_array_muxed2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_251 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_252;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_array_muxed3 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[4:0])
		1'd0: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		2'd3: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd4: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd7: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		4'd8: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		4'd9: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd10: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd11: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd12: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd13: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd14: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd15: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd16: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd17: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd18: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd19: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd20: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd21: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd22: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd23: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd24: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd25: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd26: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd27: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd28: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd29: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd30: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
		default: begin
			builder_sync_f_rhs_array_muxed3 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_252 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_253;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed1 <= 4'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[7:5])
		1'd0: begin
			builder_sync_rhs_array_muxed1 <= 3'd4;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed1 <= 4'd9;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed1 <= 3'd5;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed1 <= 2'd3;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed1 <= 2'd2;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed1 <= 4'd10;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed1 <= 3'd6;
		end
		default: begin
			builder_sync_rhs_array_muxed1 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_253 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_254;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed2 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[7:5])
		1'd0: begin
			builder_sync_rhs_array_muxed2 <= 1'd1;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed2 <= 1'd0;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed2 <= 1'd0;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed2 <= 1'd0;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed2 <= 1'd1;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed2 <= 1'd0;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed2 <= 1'd0;
		end
		default: begin
			builder_sync_rhs_array_muxed2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_254 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_255;
// synthesis translate_on
always @(*) begin
	builder_sync_f_rhs_array_muxed4 <= 1'd0;
	case (main_genericstandalone_pcs_transmitpath_d1[7:5])
		1'd0: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd1;
		end
		1'd1: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd0;
		end
		2'd2: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd0;
		end
		2'd3: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd1;
		end
		3'd4: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd1;
		end
		3'd5: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd0;
		end
		3'd6: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd0;
		end
		default: begin
			builder_sync_f_rhs_array_muxed4 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_255 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_256;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed0 <= 1'd0;
	case (main_rtio_core_outputs_channel_r0)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed0 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_256 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_257;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed1 <= 1'd0;
	case (main_rtio_core_outputs_channel_r1)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed1 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_257 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_258;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed2 <= 1'd0;
	case (main_rtio_core_outputs_channel_r2)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed2 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_258 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_259;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed3 <= 1'd0;
	case (main_rtio_core_outputs_channel_r3)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed3 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_259 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_260;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed4 <= 1'd0;
	case (main_rtio_core_outputs_channel_r4)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed4 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_260 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_261;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed5 <= 1'd0;
	case (main_rtio_core_outputs_channel_r5)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed5 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_261 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_262;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed6 <= 1'd0;
	case (main_rtio_core_outputs_channel_r6)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed6 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_262 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_263;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed7 <= 1'd0;
	case (main_rtio_core_outputs_channel_r7)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x7_inout_8x7_ointerface7_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x0_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x1_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x2_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x3_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x4_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x5_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x6_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x7_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster0_ointerface0_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x8_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x9_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x10_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x11_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x12_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster1_ointerface1_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x13_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x14_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x15_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x16_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x17_busy;
		end
		5'd28: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster2_ointerface2_busy;
		end
		5'd29: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x18_busy;
		end
		5'd30: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x19_busy;
		end
		5'd31: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x20_busy;
		end
		6'd32: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x21_busy;
		end
		6'd33: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x22_busy;
		end
		6'd34: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output0_busy;
		end
		6'd35: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output1_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed7 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_263 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_264;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed1 <= 8'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed1 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed1 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed1 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed1 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed1 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed1 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed1 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed1 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_264 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_265;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed2 <= 7'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed2 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed2 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed2 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed2 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed2 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed2 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed2 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed2 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_265 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_266;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed3 <= 8'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed3 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed3 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed3 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed3 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed3 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed3 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed3 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed3 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_266 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_267;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed4 <= 7'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed4 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed4 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed4 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed4 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed4 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed4 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed4 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed4 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_267 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_268;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed5 <= 8'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed5 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed5 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed5 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed5 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed5 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed5 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed5 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed5 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_268 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_269;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed6 <= 7'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed6 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed6 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed6 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed6 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed6 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed6 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed6 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_269 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_270;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed7 <= 8'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed7 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed7 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed7 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed7 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed7 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed7 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed7 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed7 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_270 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_271;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed8 <= 7'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed8 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed8 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed8 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed8 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed8 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed8 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed8 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed8 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_271 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_272;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed9 <= 8'd0;
	case (main_inout_8x4_inout_8x4_ointerface4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed9 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed9 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed9 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed9 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed9 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed9 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed9 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed9 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_272 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_273;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed10 <= 7'd0;
	case (main_inout_8x4_inout_8x4_ointerface4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed10 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed10 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed10 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed10 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed10 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed10 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed10 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed10 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_273 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_274;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed11 <= 8'd0;
	case (main_inout_8x5_inout_8x5_ointerface5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed11 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed11 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed11 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed11 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed11 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed11 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed11 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed11 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_274 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_275;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed12 <= 7'd0;
	case (main_inout_8x5_inout_8x5_ointerface5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed12 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed12 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed12 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed12 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed12 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed12 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed12 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_275 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_276;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed13 <= 8'd0;
	case (main_inout_8x6_inout_8x6_ointerface6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed13 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed13 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed13 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed13 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed13 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed13 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed13 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed13 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_276 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_277;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed14 <= 7'd0;
	case (main_inout_8x6_inout_8x6_ointerface6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed14 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed14 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed14 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed14 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed14 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed14 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed14 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed14 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_277 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_278;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed15 <= 8'd0;
	case (main_inout_8x7_inout_8x7_ointerface7_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed15 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed15 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed15 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed15 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed15 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed15 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed15 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed15 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_278 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_279;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed16 <= 7'd0;
	case (main_inout_8x7_inout_8x7_ointerface7_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed16 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed16 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed16 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed16 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed16 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed16 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed16 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed16 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_279 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_280;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed17 <= 8'd0;
	case (main_output_8x0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed17 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed17 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed17 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed17 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed17 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed17 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed17 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed17 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_280 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_281;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed18 <= 7'd0;
	case (main_output_8x0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed18 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed18 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed18 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed18 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed18 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed18 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed18 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed18 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_281 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_282;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed19 <= 8'd0;
	case (main_output_8x1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed19 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed19 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed19 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed19 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed19 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed19 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed19 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed19 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_282 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_283;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed20 <= 7'd0;
	case (main_output_8x1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed20 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed20 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed20 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed20 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed20 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed20 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed20 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_283 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_284;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed21 <= 8'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed21 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed21 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed21 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed21 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed21 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed21 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed21 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed21 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_284 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_285;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed22 <= 7'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed22 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed22 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed22 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed22 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed22 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed22 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed22 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed22 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_285 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_286;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed23 <= 8'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed23 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed23 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed23 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed23 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed23 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed23 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed23 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed23 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_286 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_287;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed24 <= 7'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed24 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed24 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed24 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed24 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed24 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed24 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed24 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed24 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_287 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_288;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed25 <= 8'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed25 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed25 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed25 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed25 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed25 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed25 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed25 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed25 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_288 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_289;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed26 <= 7'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed26 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed26 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed26 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed26 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed26 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed26 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed26 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_289 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_290;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed27 <= 8'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed27 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed27 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed27 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed27 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed27 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed27 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed27 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed27 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_290 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_291;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed28 <= 7'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed28 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed28 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed28 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed28 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed28 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed28 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed28 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed28 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_291 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_292;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed29 <= 8'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed29 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed29 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed29 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed29 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed29 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed29 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed29 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed29 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_292 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_293;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed30 <= 7'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed30 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed30 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed30 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed30 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed30 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed30 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed30 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed30 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_293 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_294;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed31 <= 8'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed31 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed31 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed31 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed31 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed31 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed31 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed31 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed31 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_294 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_295;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed32 <= 7'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed32 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed32 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed32 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed32 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed32 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed32 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed32 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed32 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_295 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_296;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed33 <= 8'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed33 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed33 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed33 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed33 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed33 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed33 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed33 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed33 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_296 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_297;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed34 <= 7'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed34 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed34 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed34 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed34 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed34 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed34 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed34 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed34 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_297 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_298;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed35 <= 8'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed35 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed35 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed35 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed35 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed35 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed35 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed35 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed35 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_298 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_299;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed36 <= 7'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed36 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed36 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed36 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed36 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed36 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed36 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed36 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed36 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_299 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_300;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed37 <= 8'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed37 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed37 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed37 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed37 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed37 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed37 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed37 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed37 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_300 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_301;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed38 <= 7'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed38 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed38 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed38 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed38 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed38 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed38 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed38 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed38 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_301 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_302;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed39 <= 8'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed39 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed39 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed39 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed39 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed39 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed39 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed39 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed39 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_302 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_303;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed40 <= 7'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed40 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed40 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed40 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed40 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed40 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed40 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed40 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed40 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_303 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_304;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed41 <= 8'd0;
	case (main_output_8x12_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed41 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed41 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed41 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed41 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed41 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed41 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed41 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed41 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_304 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_305;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed42 <= 7'd0;
	case (main_output_8x12_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed42 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed42 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed42 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed42 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed42 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed42 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed42 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed42 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_305 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_306;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed43 <= 8'd0;
	case (main_output_8x13_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed43 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed43 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed43 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed43 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed43 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed43 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed43 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed43 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_306 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_307;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed44 <= 7'd0;
	case (main_output_8x13_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed44 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed44 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed44 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed44 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed44 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed44 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed44 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed44 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_307 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_308;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed45 <= 8'd0;
	case (main_output_8x14_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed45 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed45 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed45 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed45 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed45 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed45 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed45 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed45 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_308 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_309;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed46 <= 7'd0;
	case (main_output_8x14_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed46 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed46 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed46 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed46 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed46 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed46 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed46 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed46 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_309 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_310;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed47 <= 8'd0;
	case (main_output_8x15_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed47 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed47 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed47 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed47 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed47 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed47 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed47 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed47 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_310 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_311;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed48 <= 7'd0;
	case (main_output_8x15_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed48 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed48 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed48 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed48 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed48 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed48 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed48 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed48 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_311 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_312;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed49 <= 8'd0;
	case (main_output_8x16_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed49 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed49 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed49 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed49 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed49 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed49 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed49 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed49 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_312 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_313;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed50 <= 7'd0;
	case (main_output_8x16_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed50 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed50 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed50 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed50 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed50 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed50 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed50 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed50 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_313 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_314;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed51 <= 8'd0;
	case (main_output_8x17_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed51 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed51 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed51 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed51 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed51 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed51 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed51 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed51 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_314 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_315;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed52 <= 7'd0;
	case (main_output_8x17_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed52 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed52 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed52 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed52 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed52 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed52 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed52 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed52 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_315 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_316;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed53 <= 8'd0;
	case (main_output_8x18_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed53 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed53 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed53 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed53 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed53 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed53 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed53 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed53 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_316 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_317;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed54 <= 7'd0;
	case (main_output_8x18_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed54 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed54 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed54 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed54 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed54 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed54 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed54 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed54 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_317 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_318;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed55 <= 8'd0;
	case (main_output_8x19_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed55 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed55 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed55 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed55 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed55 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed55 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed55 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed55 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_318 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_319;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed56 <= 7'd0;
	case (main_output_8x19_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed56 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed56 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed56 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed56 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed56 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed56 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed56 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed56 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_319 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_320;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed57 <= 8'd0;
	case (main_output_8x20_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed57 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed57 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed57 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed57 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed57 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed57 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed57 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed57 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_320 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_321;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed58 <= 7'd0;
	case (main_output_8x20_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed58 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed58 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed58 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed58 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed58 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed58 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed58 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed58 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_321 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_322;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed59 <= 8'd0;
	case (main_output_8x21_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed59 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed59 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed59 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed59 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed59 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed59 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed59 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed59 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_322 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_323;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed60 <= 7'd0;
	case (main_output_8x21_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed60 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed60 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed60 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed60 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed60 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed60 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed60 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed60 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_323 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_324;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed61 <= 8'd0;
	case (main_output_8x22_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed61 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed61 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed61 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed61 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed61 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed61 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed61 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed61 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_324 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_325;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed62 <= 7'd0;
	case (main_output_8x22_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed62 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed62 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed62 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed62 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed62 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed62 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed62 <= 6'd63;
		end
		default: begin
			builder_sync_f_t_array_muxed62 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_325 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_326;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed3 <= 61'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			builder_sync_rhs_array_muxed3 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_326 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_327;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed4 <= 61'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane_plus_one)
		1'd0: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			builder_sync_rhs_array_muxed4 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_327 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_328;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed1 <= 32'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record0_fifo_out_data;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record1_fifo_out_data;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record2_fifo_out_data;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record3_fifo_out_data;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record4_fifo_out_data;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record5_fifo_out_data;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record6_fifo_out_data;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record7_fifo_out_data;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record8_fifo_out_data;
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record9_fifo_out_data;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_array_muxed1 <= main_rtio_core_inputs_record10_fifo_out_data;
		end
		5'd29: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd31: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd32: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd33: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd34: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd35: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_328 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_329;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed2 <= 65'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record0_fifo_out_timestamp <<< 1'd0);
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record1_fifo_out_timestamp <<< 1'd0);
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record2_fifo_out_timestamp <<< 1'd0);
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record3_fifo_out_timestamp <<< 1'd0);
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record4_fifo_out_timestamp <<< 1'd0);
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record5_fifo_out_timestamp <<< 1'd0);
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record6_fifo_out_timestamp <<< 1'd0);
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed2 <= (main_rtio_core_inputs_record7_fifo_out_timestamp <<< 1'd0);
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd28: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd29: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd30: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd31: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd32: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd33: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd34: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd35: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed2 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_329 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_330;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed5 <= 32'd0;
	case (main_genericstandalone_mailbox_i1_adr[1:0])
		1'd0: begin
			builder_sync_rhs_array_muxed5 <= main_genericstandalone_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed5 <= main_genericstandalone_mailbox1;
		end
		default: begin
			builder_sync_rhs_array_muxed5 <= main_genericstandalone_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_330 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_331;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed6 <= 32'd0;
	case (main_genericstandalone_mailbox_i2_adr[1:0])
		1'd0: begin
			builder_sync_rhs_array_muxed6 <= main_genericstandalone_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed6 <= main_genericstandalone_mailbox1;
		end
		default: begin
			builder_sync_rhs_array_muxed6 <= main_genericstandalone_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_331 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_332;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed4 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed4 <= main_mon_bussynchronizer0_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed4 <= main_mon_bussynchronizer1_o;
		end
	endcase
// synthesis translate_off
	dummy_d_332 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_333;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed5 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed5 <= main_mon_bussynchronizer2_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed5 <= main_mon_bussynchronizer3_o;
		end
	endcase
// synthesis translate_off
	dummy_d_333 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_334;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed6 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed6 <= main_mon_bussynchronizer4_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed6 <= main_mon_bussynchronizer5_o;
		end
	endcase
// synthesis translate_off
	dummy_d_334 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_335;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed7 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed7 <= main_mon_bussynchronizer6_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed7 <= main_mon_bussynchronizer7_o;
		end
	endcase
// synthesis translate_off
	dummy_d_335 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_336;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed8 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed8 <= main_mon_bussynchronizer8_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed8 <= main_mon_bussynchronizer9_o;
		end
	endcase
// synthesis translate_off
	dummy_d_336 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_337;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed9 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed9 <= main_mon_bussynchronizer10_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed9 <= main_mon_bussynchronizer11_o;
		end
	endcase
// synthesis translate_off
	dummy_d_337 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_338;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed10 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed10 <= main_mon_bussynchronizer12_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed10 <= main_mon_bussynchronizer13_o;
		end
	endcase
// synthesis translate_off
	dummy_d_338 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_339;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed11 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed11 <= main_mon_bussynchronizer14_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed11 <= main_mon_bussynchronizer15_o;
		end
	endcase
// synthesis translate_off
	dummy_d_339 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_340;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed12 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed12 <= main_mon_bussynchronizer16_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_340 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_341;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed13 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed13 <= main_mon_bussynchronizer17_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_341 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_342;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed14 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed14 <= main_mon_bussynchronizer18_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_342 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_343;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed15 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed15 <= main_mon_bussynchronizer19_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_343 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_344;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed16 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed16 <= main_mon_bussynchronizer20_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_344 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_345;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed17 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed17 <= main_mon_bussynchronizer21_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_345 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_346;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed18 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed18 <= main_mon_bussynchronizer22_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_346 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_347;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed19 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed19 <= main_mon_bussynchronizer23_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_347 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_348;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed20 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_348 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_349;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed21 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed21 <= main_mon_bussynchronizer24_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_349 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_350;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed22 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed22 <= main_mon_bussynchronizer25_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_350 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_351;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed23 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed23 <= main_mon_bussynchronizer26_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_351 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_352;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed24 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed24 <= main_mon_bussynchronizer27_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_352 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_353;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed25 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed25 <= main_mon_bussynchronizer28_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_353 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_354;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed26 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_354 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_355;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed27 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed27 <= main_mon_bussynchronizer29_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_355 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_356;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed28 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed28 <= main_mon_bussynchronizer30_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_356 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_357;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed29 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed29 <= main_mon_bussynchronizer31_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_357 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_358;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed30 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer32_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_358 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_359;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed31 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed31 <= main_mon_bussynchronizer33_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_359 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_360;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed32 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed32 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_360 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_361;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed33 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed33 <= main_mon_bussynchronizer34_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_361 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_362;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed34 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed34 <= main_mon_bussynchronizer35_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_362 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_363;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed35 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed35 <= main_mon_bussynchronizer36_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed35 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_363 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_364;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed36 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed36 <= main_mon_bussynchronizer37_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_364 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_365;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed37 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed37 <= main_mon_bussynchronizer38_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_365 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_366;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed38 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed38 <= main_mon_bussynchronizer39_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_366 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_367;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed39 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed39 <= main_mon_bussynchronizer40_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_367 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_368;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed40 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed40 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_368 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_369;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed3 <= 1'd0;
	case (main_mon_chan_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed4;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed5;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed6;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed7;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed8;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed9;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed10;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed11;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed12;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed13;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed14;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed15;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed16;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed17;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed18;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed19;
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed20;
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed21;
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed22;
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed23;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed24;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed25;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed26;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed27;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed28;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed29;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed30;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed31;
		end
		5'd28: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed32;
		end
		5'd29: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed33;
		end
		5'd30: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed34;
		end
		5'd31: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed35;
		end
		6'd32: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed36;
		end
		6'd33: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed37;
		end
		6'd34: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed38;
		end
		6'd35: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed39;
		end
		default: begin
			builder_sync_t_rhs_array_muxed3 <= builder_sync_t_rhs_array_muxed40;
		end
	endcase
// synthesis translate_off
	dummy_d_369 <= dummy_s;
// synthesis translate_on
end
assign main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx = builder_xilinxmultiregimpl0_regs1;
assign builder_xilinxasyncresetsynchronizerimpl0 = (~main_genericstandalone_genericstandalone_pll_locked);
assign main_genericstandalone_pcs_seen_valid_ci_toggle_o = builder_xilinxmultiregimpl1_regs1;
assign main_genericstandalone_pcs_rx_config_reg_toggle_o = builder_xilinxmultiregimpl2_regs1;
assign main_genericstandalone_pcs_rx_config_reg_ack_toggle_o = builder_xilinxmultiregimpl3_regs1;
assign builder_xilinxasyncresetsynchronizerimpl1 = (~main_genericstandalone_tx_mmcm_locked);
assign builder_xilinxasyncresetsynchronizerimpl2 = (~main_genericstandalone_rx_mmcm_locked);
assign main_genericstandalone_tx_init_qpll_lock1 = builder_xilinxmultiregimpl4_regs1;
assign main_genericstandalone_rx_init_rx_pma_reset_done1 = builder_xilinxmultiregimpl5_regs1;
assign main_genericstandalone_toggle_o = builder_xilinxmultiregimpl6_regs1;
assign main_genericstandalone_ps_preamble_error_toggle_o = builder_xilinxmultiregimpl7_regs1;
assign main_genericstandalone_ps_crc_error_toggle_o = builder_xilinxmultiregimpl8_regs1;
assign main_genericstandalone_tx_cdc_produce_rdomain = builder_xilinxmultiregimpl9_regs1;
assign main_genericstandalone_tx_cdc_consume_wdomain = builder_xilinxmultiregimpl10_regs1;
assign main_genericstandalone_rx_cdc_produce_rdomain = builder_xilinxmultiregimpl11_regs1;
assign main_genericstandalone_rx_cdc_consume_wdomain = builder_xilinxmultiregimpl12_regs1;
assign main_i2c_status1 = builder_xilinxmultiregimpl13_regs1;
assign main_i2c_status2 = builder_xilinxmultiregimpl14_regs1;
assign builder_xilinxasyncresetsynchronizerimpl3 = (~main_rtio_crg_pll_locked);
assign main_rtio_crg_pll_locked_status = builder_xilinxmultiregimpl15_regs1;
assign main_rtio_tsc_value_gray_sys = builder_xilinxmultiregimpl16_regs1;
assign main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain = builder_xilinxmultiregimpl17_regs1;
assign main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain = builder_xilinxmultiregimpl18_regs1;
assign main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain = builder_xilinxmultiregimpl19_regs1;
assign main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain = builder_xilinxmultiregimpl20_regs1;
assign main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain = builder_xilinxmultiregimpl21_regs1;
assign main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain = builder_xilinxmultiregimpl22_regs1;
assign main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain = builder_xilinxmultiregimpl23_regs1;
assign main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain = builder_xilinxmultiregimpl24_regs1;
assign main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain = builder_xilinxmultiregimpl25_regs1;
assign main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain = builder_xilinxmultiregimpl26_regs1;
assign main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain = builder_xilinxmultiregimpl27_regs1;
assign main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain = builder_xilinxmultiregimpl28_regs1;
assign main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain = builder_xilinxmultiregimpl29_regs1;
assign main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain = builder_xilinxmultiregimpl30_regs1;
assign main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain = builder_xilinxmultiregimpl31_regs1;
assign main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain = builder_xilinxmultiregimpl32_regs1;
assign main_rtio_core_inputs_asyncfifo0_produce_rdomain = builder_xilinxmultiregimpl33_regs1;
assign main_rtio_core_inputs_asyncfifo0_consume_wdomain = builder_xilinxmultiregimpl34_regs1;
assign main_rtio_core_inputs_blindtransfer0_ps_toggle_o = builder_xilinxmultiregimpl35_regs1;
assign main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o = builder_xilinxmultiregimpl36_regs1;
assign main_rtio_core_inputs_asyncfifo1_produce_rdomain = builder_xilinxmultiregimpl37_regs1;
assign main_rtio_core_inputs_asyncfifo1_consume_wdomain = builder_xilinxmultiregimpl38_regs1;
assign main_rtio_core_inputs_blindtransfer1_ps_toggle_o = builder_xilinxmultiregimpl39_regs1;
assign main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o = builder_xilinxmultiregimpl40_regs1;
assign main_rtio_core_inputs_asyncfifo2_produce_rdomain = builder_xilinxmultiregimpl41_regs1;
assign main_rtio_core_inputs_asyncfifo2_consume_wdomain = builder_xilinxmultiregimpl42_regs1;
assign main_rtio_core_inputs_blindtransfer2_ps_toggle_o = builder_xilinxmultiregimpl43_regs1;
assign main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o = builder_xilinxmultiregimpl44_regs1;
assign main_rtio_core_inputs_asyncfifo3_produce_rdomain = builder_xilinxmultiregimpl45_regs1;
assign main_rtio_core_inputs_asyncfifo3_consume_wdomain = builder_xilinxmultiregimpl46_regs1;
assign main_rtio_core_inputs_blindtransfer3_ps_toggle_o = builder_xilinxmultiregimpl47_regs1;
assign main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o = builder_xilinxmultiregimpl48_regs1;
assign main_rtio_core_inputs_asyncfifo4_produce_rdomain = builder_xilinxmultiregimpl49_regs1;
assign main_rtio_core_inputs_asyncfifo4_consume_wdomain = builder_xilinxmultiregimpl50_regs1;
assign main_rtio_core_inputs_blindtransfer4_ps_toggle_o = builder_xilinxmultiregimpl51_regs1;
assign main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o = builder_xilinxmultiregimpl52_regs1;
assign main_rtio_core_inputs_asyncfifo5_produce_rdomain = builder_xilinxmultiregimpl53_regs1;
assign main_rtio_core_inputs_asyncfifo5_consume_wdomain = builder_xilinxmultiregimpl54_regs1;
assign main_rtio_core_inputs_blindtransfer5_ps_toggle_o = builder_xilinxmultiregimpl55_regs1;
assign main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o = builder_xilinxmultiregimpl56_regs1;
assign main_rtio_core_inputs_asyncfifo6_produce_rdomain = builder_xilinxmultiregimpl57_regs1;
assign main_rtio_core_inputs_asyncfifo6_consume_wdomain = builder_xilinxmultiregimpl58_regs1;
assign main_rtio_core_inputs_blindtransfer6_ps_toggle_o = builder_xilinxmultiregimpl59_regs1;
assign main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o = builder_xilinxmultiregimpl60_regs1;
assign main_rtio_core_inputs_asyncfifo7_produce_rdomain = builder_xilinxmultiregimpl61_regs1;
assign main_rtio_core_inputs_asyncfifo7_consume_wdomain = builder_xilinxmultiregimpl62_regs1;
assign main_rtio_core_inputs_blindtransfer7_ps_toggle_o = builder_xilinxmultiregimpl63_regs1;
assign main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o = builder_xilinxmultiregimpl64_regs1;
assign main_rtio_core_inputs_asyncfifo8_produce_rdomain = builder_xilinxmultiregimpl65_regs1;
assign main_rtio_core_inputs_asyncfifo8_consume_wdomain = builder_xilinxmultiregimpl66_regs1;
assign main_rtio_core_inputs_blindtransfer8_ps_toggle_o = builder_xilinxmultiregimpl67_regs1;
assign main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o = builder_xilinxmultiregimpl68_regs1;
assign main_rtio_core_inputs_asyncfifo9_produce_rdomain = builder_xilinxmultiregimpl69_regs1;
assign main_rtio_core_inputs_asyncfifo9_consume_wdomain = builder_xilinxmultiregimpl70_regs1;
assign main_rtio_core_inputs_blindtransfer9_ps_toggle_o = builder_xilinxmultiregimpl71_regs1;
assign main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o = builder_xilinxmultiregimpl72_regs1;
assign main_rtio_core_inputs_asyncfifo10_produce_rdomain = builder_xilinxmultiregimpl73_regs1;
assign main_rtio_core_inputs_asyncfifo10_consume_wdomain = builder_xilinxmultiregimpl74_regs1;
assign main_rtio_core_inputs_blindtransfer10_ps_toggle_o = builder_xilinxmultiregimpl75_regs1;
assign main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o = builder_xilinxmultiregimpl76_regs1;
assign main_rtio_core_o_collision_sync_ps_toggle_o = builder_xilinxmultiregimpl77_regs1;
assign main_rtio_core_o_collision_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl78_regs1;
assign main_rtio_core_o_collision_sync_data_o = builder_xilinxmultiregimpl79_regs1;
assign main_rtio_core_o_busy_sync_ps_toggle_o = builder_xilinxmultiregimpl80_regs1;
assign main_rtio_core_o_busy_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl81_regs1;
assign main_rtio_core_o_busy_sync_data_o = builder_xilinxmultiregimpl82_regs1;
assign main_mon_bussynchronizer0_o = builder_xilinxmultiregimpl83_regs1;
assign main_mon_bussynchronizer1_o = builder_xilinxmultiregimpl84_regs1;
assign main_mon_bussynchronizer2_o = builder_xilinxmultiregimpl85_regs1;
assign main_mon_bussynchronizer3_o = builder_xilinxmultiregimpl86_regs1;
assign main_mon_bussynchronizer4_o = builder_xilinxmultiregimpl87_regs1;
assign main_mon_bussynchronizer5_o = builder_xilinxmultiregimpl88_regs1;
assign main_mon_bussynchronizer6_o = builder_xilinxmultiregimpl89_regs1;
assign main_mon_bussynchronizer7_o = builder_xilinxmultiregimpl90_regs1;
assign main_mon_bussynchronizer8_o = builder_xilinxmultiregimpl91_regs1;
assign main_mon_bussynchronizer9_o = builder_xilinxmultiregimpl92_regs1;
assign main_mon_bussynchronizer10_o = builder_xilinxmultiregimpl93_regs1;
assign main_mon_bussynchronizer11_o = builder_xilinxmultiregimpl94_regs1;
assign main_mon_bussynchronizer12_o = builder_xilinxmultiregimpl95_regs1;
assign main_mon_bussynchronizer13_o = builder_xilinxmultiregimpl96_regs1;
assign main_mon_bussynchronizer14_o = builder_xilinxmultiregimpl97_regs1;
assign main_mon_bussynchronizer15_o = builder_xilinxmultiregimpl98_regs1;
assign main_mon_bussynchronizer16_o = builder_xilinxmultiregimpl99_regs1;
assign main_mon_bussynchronizer17_o = builder_xilinxmultiregimpl100_regs1;
assign main_mon_bussynchronizer18_o = builder_xilinxmultiregimpl101_regs1;
assign main_mon_bussynchronizer19_o = builder_xilinxmultiregimpl102_regs1;
assign main_mon_bussynchronizer20_o = builder_xilinxmultiregimpl103_regs1;
assign main_mon_bussynchronizer21_o = builder_xilinxmultiregimpl104_regs1;
assign main_mon_bussynchronizer22_o = builder_xilinxmultiregimpl105_regs1;
assign main_mon_bussynchronizer23_o = builder_xilinxmultiregimpl106_regs1;
assign main_mon_bussynchronizer24_o = builder_xilinxmultiregimpl107_regs1;
assign main_mon_bussynchronizer25_o = builder_xilinxmultiregimpl108_regs1;
assign main_mon_bussynchronizer26_o = builder_xilinxmultiregimpl109_regs1;
assign main_mon_bussynchronizer27_o = builder_xilinxmultiregimpl110_regs1;
assign main_mon_bussynchronizer28_o = builder_xilinxmultiregimpl111_regs1;
assign main_mon_bussynchronizer29_o = builder_xilinxmultiregimpl112_regs1;
assign main_mon_bussynchronizer30_o = builder_xilinxmultiregimpl113_regs1;
assign main_mon_bussynchronizer31_o = builder_xilinxmultiregimpl114_regs1;
assign main_mon_bussynchronizer32_o = builder_xilinxmultiregimpl115_regs1;
assign main_mon_bussynchronizer33_o = builder_xilinxmultiregimpl116_regs1;
assign main_mon_bussynchronizer34_o = builder_xilinxmultiregimpl117_regs1;
assign main_mon_bussynchronizer35_o = builder_xilinxmultiregimpl118_regs1;
assign main_mon_bussynchronizer36_o = builder_xilinxmultiregimpl119_regs1;
assign main_mon_bussynchronizer37_o = builder_xilinxmultiregimpl120_regs1;
assign main_mon_bussynchronizer38_o = builder_xilinxmultiregimpl121_regs1;
assign main_mon_bussynchronizer39_o = builder_xilinxmultiregimpl122_regs1;
assign main_mon_bussynchronizer40_o = builder_xilinxmultiregimpl123_regs1;
assign main_inout_8x0_inout_8x0_override_en = builder_xilinxmultiregimpl124_regs1;
assign main_inout_8x0_inout_8x0_override_o = builder_xilinxmultiregimpl125_regs1;
assign main_inout_8x0_inout_8x0_override_oe = builder_xilinxmultiregimpl126_regs1;
assign main_inout_8x1_inout_8x1_override_en = builder_xilinxmultiregimpl127_regs1;
assign main_inout_8x1_inout_8x1_override_o = builder_xilinxmultiregimpl128_regs1;
assign main_inout_8x1_inout_8x1_override_oe = builder_xilinxmultiregimpl129_regs1;
assign main_inout_8x2_inout_8x2_override_en = builder_xilinxmultiregimpl130_regs1;
assign main_inout_8x2_inout_8x2_override_o = builder_xilinxmultiregimpl131_regs1;
assign main_inout_8x2_inout_8x2_override_oe = builder_xilinxmultiregimpl132_regs1;
assign main_inout_8x3_inout_8x3_override_en = builder_xilinxmultiregimpl133_regs1;
assign main_inout_8x3_inout_8x3_override_o = builder_xilinxmultiregimpl134_regs1;
assign main_inout_8x3_inout_8x3_override_oe = builder_xilinxmultiregimpl135_regs1;
assign main_inout_8x4_inout_8x4_override_en = builder_xilinxmultiregimpl136_regs1;
assign main_inout_8x4_inout_8x4_override_o = builder_xilinxmultiregimpl137_regs1;
assign main_inout_8x4_inout_8x4_override_oe = builder_xilinxmultiregimpl138_regs1;
assign main_inout_8x5_inout_8x5_override_en = builder_xilinxmultiregimpl139_regs1;
assign main_inout_8x5_inout_8x5_override_o = builder_xilinxmultiregimpl140_regs1;
assign main_inout_8x5_inout_8x5_override_oe = builder_xilinxmultiregimpl141_regs1;
assign main_inout_8x6_inout_8x6_override_en = builder_xilinxmultiregimpl142_regs1;
assign main_inout_8x6_inout_8x6_override_o = builder_xilinxmultiregimpl143_regs1;
assign main_inout_8x6_inout_8x6_override_oe = builder_xilinxmultiregimpl144_regs1;
assign main_inout_8x7_inout_8x7_override_en = builder_xilinxmultiregimpl145_regs1;
assign main_inout_8x7_inout_8x7_override_o = builder_xilinxmultiregimpl146_regs1;
assign main_inout_8x7_inout_8x7_override_oe = builder_xilinxmultiregimpl147_regs1;
assign main_output_8x0_override_en = builder_xilinxmultiregimpl148_regs1;
assign main_output_8x0_override_o = builder_xilinxmultiregimpl149_regs1;
assign main_output_8x1_override_en = builder_xilinxmultiregimpl150_regs1;
assign main_output_8x1_override_o = builder_xilinxmultiregimpl151_regs1;
assign main_output_8x2_override_en = builder_xilinxmultiregimpl152_regs1;
assign main_output_8x2_override_o = builder_xilinxmultiregimpl153_regs1;
assign main_output_8x3_override_en = builder_xilinxmultiregimpl154_regs1;
assign main_output_8x3_override_o = builder_xilinxmultiregimpl155_regs1;
assign main_output_8x4_override_en = builder_xilinxmultiregimpl156_regs1;
assign main_output_8x4_override_o = builder_xilinxmultiregimpl157_regs1;
assign main_output_8x5_override_en = builder_xilinxmultiregimpl158_regs1;
assign main_output_8x5_override_o = builder_xilinxmultiregimpl159_regs1;
assign main_output_8x6_override_en = builder_xilinxmultiregimpl160_regs1;
assign main_output_8x6_override_o = builder_xilinxmultiregimpl161_regs1;
assign main_output_8x7_override_en = builder_xilinxmultiregimpl162_regs1;
assign main_output_8x7_override_o = builder_xilinxmultiregimpl163_regs1;
assign main_output_8x8_override_en = builder_xilinxmultiregimpl164_regs1;
assign main_output_8x8_override_o = builder_xilinxmultiregimpl165_regs1;
assign main_output_8x9_override_en = builder_xilinxmultiregimpl166_regs1;
assign main_output_8x9_override_o = builder_xilinxmultiregimpl167_regs1;
assign main_output_8x10_override_en = builder_xilinxmultiregimpl168_regs1;
assign main_output_8x10_override_o = builder_xilinxmultiregimpl169_regs1;
assign main_output_8x11_override_en = builder_xilinxmultiregimpl170_regs1;
assign main_output_8x11_override_o = builder_xilinxmultiregimpl171_regs1;
assign main_output_8x12_override_en = builder_xilinxmultiregimpl172_regs1;
assign main_output_8x12_override_o = builder_xilinxmultiregimpl173_regs1;
assign main_output_8x13_override_en = builder_xilinxmultiregimpl174_regs1;
assign main_output_8x13_override_o = builder_xilinxmultiregimpl175_regs1;
assign main_output_8x14_override_en = builder_xilinxmultiregimpl176_regs1;
assign main_output_8x14_override_o = builder_xilinxmultiregimpl177_regs1;
assign main_output_8x15_override_en = builder_xilinxmultiregimpl178_regs1;
assign main_output_8x15_override_o = builder_xilinxmultiregimpl179_regs1;
assign main_output_8x16_override_en = builder_xilinxmultiregimpl180_regs1;
assign main_output_8x16_override_o = builder_xilinxmultiregimpl181_regs1;
assign main_output_8x17_override_en = builder_xilinxmultiregimpl182_regs1;
assign main_output_8x17_override_o = builder_xilinxmultiregimpl183_regs1;
assign main_output_8x18_override_en = builder_xilinxmultiregimpl184_regs1;
assign main_output_8x18_override_o = builder_xilinxmultiregimpl185_regs1;
assign main_output_8x19_override_en = builder_xilinxmultiregimpl186_regs1;
assign main_output_8x19_override_o = builder_xilinxmultiregimpl187_regs1;
assign main_output_8x20_override_en = builder_xilinxmultiregimpl188_regs1;
assign main_output_8x20_override_o = builder_xilinxmultiregimpl189_regs1;
assign main_output_8x21_override_en = builder_xilinxmultiregimpl190_regs1;
assign main_output_8x21_override_o = builder_xilinxmultiregimpl191_regs1;
assign main_output_8x22_override_en = builder_xilinxmultiregimpl192_regs1;
assign main_output_8x22_override_o = builder_xilinxmultiregimpl193_regs1;
assign main_output0_override_en = builder_xilinxmultiregimpl194_regs1;
assign main_output0_override_o = builder_xilinxmultiregimpl195_regs1;
assign main_output1_override_en = builder_xilinxmultiregimpl196_regs1;
assign main_output1_override_o = builder_xilinxmultiregimpl197_regs1;

always @(posedge clk200_clk) begin
	if ((main_genericstandalone_genericstandalone_reset_counter != 1'd0)) begin
		main_genericstandalone_genericstandalone_reset_counter <= (main_genericstandalone_genericstandalone_reset_counter - 1'd1);
	end else begin
		main_genericstandalone_genericstandalone_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		main_genericstandalone_genericstandalone_reset_counter <= 4'd15;
		main_genericstandalone_genericstandalone_ic_reset <= 1'd1;
	end
end

always @(posedge eth_rx_clk) begin
	main_genericstandalone_pcs_rx_en_d <= main_genericstandalone_pcs_receivepath_rx_en;
	main_genericstandalone_pcs_source_stb <= main_genericstandalone_pcs_receivepath_rx_en;
	main_genericstandalone_pcs_source_payload_data <= main_genericstandalone_pcs_receivepath_rx_data;
	if (main_genericstandalone_pcs_receivepath_seen_config_reg) begin
		main_genericstandalone_pcs_c_counter <= 3'd4;
	end else begin
		if ((main_genericstandalone_pcs_c_counter != 1'd0)) begin
			main_genericstandalone_pcs_c_counter <= (main_genericstandalone_pcs_c_counter - 1'd1);
		end
	end
	main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd0;
	main_genericstandalone_pcs_rx_config_reg_i <= 1'd0;
	if (main_genericstandalone_pcs_receivepath_seen_config_reg) begin
		main_genericstandalone_pcs_previous_config_reg <= main_genericstandalone_pcs_receivepath_config_reg;
		if (((main_genericstandalone_pcs_c_counter == 1'd1) & (main_genericstandalone_pcs_previous_config_reg == main_genericstandalone_pcs_receivepath_config_reg))) begin
			if (main_genericstandalone_pcs_previous_config_reg[14]) begin
				main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd1;
			end else begin
				main_genericstandalone_pcs_rx_config_reg_i <= 1'd1;
			end
		end
	end
	main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd0;
	if (main_genericstandalone_pcs_receivepath_load_config_reg_lsb) begin
		main_genericstandalone_pcs_receivepath_config_reg_lsb <= main_genericstandalone_pcs_receivepath_d;
	end
	if (main_genericstandalone_pcs_receivepath_load_config_reg_msb) begin
		main_genericstandalone_pcs_receivepath_config_reg <= {main_genericstandalone_pcs_receivepath_d, main_genericstandalone_pcs_receivepath_config_reg_lsb};
		main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd1;
	end
	main_genericstandalone_pcs_receivepath_k <= 1'd0;
	if ((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] == 4'd15)) begin
		main_genericstandalone_pcs_receivepath_k <= 1'd1;
		main_genericstandalone_pcs_receivepath_code3b <= builder_sync_t_rhs_array_muxed0;
	end else begin
		if ((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] == 6'd48)) begin
			main_genericstandalone_pcs_receivepath_k <= 1'd1;
			main_genericstandalone_pcs_receivepath_code3b <= builder_sync_f_t_array_muxed0;
		end else begin
			if (((main_genericstandalone_pcs_receivepath_input_msb_first[3:0] == 3'd7) | (main_genericstandalone_pcs_receivepath_input_msb_first[3:0] == 4'd8))) begin
				if (((((((main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd35) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 5'd19)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 4'd11)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd52)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 6'd44)) & (main_genericstandalone_pcs_receivepath_input_msb_first[9:4] != 5'd28))) begin
					main_genericstandalone_pcs_receivepath_k <= 1'd1;
				end
			end
			main_genericstandalone_pcs_receivepath_code3b <= builder_sync_f_rhs_array_muxed0;
		end
	end
	main_genericstandalone_pcs_receivepath_code5b <= builder_sync_rhs_array_muxed0;
	builder_a7_1000basex_receivepath_state <= builder_a7_1000basex_receivepath_next_state;
	if (main_genericstandalone_pcs_seen_valid_ci_i) begin
		main_genericstandalone_pcs_seen_valid_ci_toggle_i <= (~main_genericstandalone_pcs_seen_valid_ci_toggle_i);
	end
	if (main_genericstandalone_pcs_rx_config_reg_i) begin
		main_genericstandalone_pcs_rx_config_reg_toggle_i <= (~main_genericstandalone_pcs_rx_config_reg_toggle_i);
	end
	if (main_genericstandalone_pcs_rx_config_reg_ack_i) begin
		main_genericstandalone_pcs_rx_config_reg_ack_toggle_i <= (~main_genericstandalone_pcs_rx_config_reg_ack_toggle_i);
	end
	if ((main_genericstandalone_phase_half == main_genericstandalone_phase_half_rereg)) begin
		main_genericstandalone_rx_data1 <= main_genericstandalone_rx_data_half[19:10];
	end else begin
		main_genericstandalone_rx_data1 <= main_genericstandalone_rx_data_half[9:0];
	end
	main_genericstandalone_phase_half <= (~main_genericstandalone_phase_half);
	builder_liteethmacpreamblechecker_state <= builder_liteethmacpreamblechecker_next_state;
	if (main_genericstandalone_crc32_checker_crc_ce) begin
		main_genericstandalone_crc32_checker_crc_reg <= main_genericstandalone_crc32_checker_crc_next;
	end
	if (main_genericstandalone_crc32_checker_crc_reset) begin
		main_genericstandalone_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable) & (~main_genericstandalone_crc32_checker_syncfifo_replace))) begin
		if ((main_genericstandalone_crc32_checker_syncfifo_produce == 3'd4)) begin
			main_genericstandalone_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			main_genericstandalone_crc32_checker_syncfifo_produce <= (main_genericstandalone_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (main_genericstandalone_crc32_checker_syncfifo_do_read) begin
		if ((main_genericstandalone_crc32_checker_syncfifo_consume == 3'd4)) begin
			main_genericstandalone_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			main_genericstandalone_crc32_checker_syncfifo_consume <= (main_genericstandalone_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((main_genericstandalone_crc32_checker_syncfifo_syncfifo_we & main_genericstandalone_crc32_checker_syncfifo_syncfifo_writable) & (~main_genericstandalone_crc32_checker_syncfifo_replace))) begin
		if ((~main_genericstandalone_crc32_checker_syncfifo_do_read)) begin
			main_genericstandalone_crc32_checker_syncfifo_level <= (main_genericstandalone_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_crc32_checker_syncfifo_do_read) begin
			main_genericstandalone_crc32_checker_syncfifo_level <= (main_genericstandalone_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (main_genericstandalone_crc32_checker_fifo_reset) begin
		main_genericstandalone_crc32_checker_syncfifo_level <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_produce <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_consume <= 3'd0;
	end
	builder_liteethmaccrc32checker_state <= builder_liteethmaccrc32checker_next_state;
	if (main_genericstandalone_ps_preamble_error_i) begin
		main_genericstandalone_ps_preamble_error_toggle_i <= (~main_genericstandalone_ps_preamble_error_toggle_i);
	end
	if (main_genericstandalone_ps_crc_error_i) begin
		main_genericstandalone_ps_crc_error_toggle_i <= (~main_genericstandalone_ps_crc_error_toggle_i);
	end
	if (main_genericstandalone_rx_converter_converter_source_ack) begin
		main_genericstandalone_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (main_genericstandalone_rx_converter_converter_load_part) begin
		if (((main_genericstandalone_rx_converter_converter_demux == 2'd3) | main_genericstandalone_rx_converter_converter_sink_eop)) begin
			main_genericstandalone_rx_converter_converter_demux <= 1'd0;
			main_genericstandalone_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			main_genericstandalone_rx_converter_converter_demux <= (main_genericstandalone_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((main_genericstandalone_rx_converter_converter_source_stb & main_genericstandalone_rx_converter_converter_source_ack)) begin
		main_genericstandalone_rx_converter_converter_source_eop <= main_genericstandalone_rx_converter_converter_sink_eop;
	end else begin
		if ((main_genericstandalone_rx_converter_converter_sink_stb & main_genericstandalone_rx_converter_converter_sink_ack)) begin
			main_genericstandalone_rx_converter_converter_source_eop <= (main_genericstandalone_rx_converter_converter_sink_eop | main_genericstandalone_rx_converter_converter_source_eop);
		end
	end
	if (main_genericstandalone_rx_converter_converter_load_part) begin
		case (main_genericstandalone_rx_converter_converter_demux)
			1'd0: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[39:30] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[29:20] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[19:10] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				main_genericstandalone_rx_converter_converter_source_payload_data[9:0] <= main_genericstandalone_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	main_genericstandalone_rx_cdc_graycounter0_q_binary <= main_genericstandalone_rx_cdc_graycounter0_q_next_binary;
	main_genericstandalone_rx_cdc_graycounter0_q <= main_genericstandalone_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		main_genericstandalone_pcs_receivepath_seen_config_reg <= 1'd0;
		main_genericstandalone_pcs_receivepath_config_reg <= 16'd0;
		main_genericstandalone_pcs_receivepath_k <= 1'd0;
		main_genericstandalone_pcs_receivepath_code5b <= 5'd0;
		main_genericstandalone_pcs_receivepath_code3b <= 3'd0;
		main_genericstandalone_pcs_receivepath_config_reg_lsb <= 8'd0;
		main_genericstandalone_pcs_source_stb <= 1'd0;
		main_genericstandalone_pcs_source_payload_data <= 8'd0;
		main_genericstandalone_pcs_rx_en_d <= 1'd0;
		main_genericstandalone_pcs_rx_config_reg_i <= 1'd0;
		main_genericstandalone_pcs_rx_config_reg_ack_i <= 1'd0;
		main_genericstandalone_pcs_c_counter <= 3'd0;
		main_genericstandalone_pcs_previous_config_reg <= 16'd0;
		main_genericstandalone_rx_data1 <= 10'd0;
		main_genericstandalone_phase_half <= 1'd0;
		main_genericstandalone_crc32_checker_crc_reg <= 32'd4294967295;
		main_genericstandalone_crc32_checker_syncfifo_level <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_produce <= 3'd0;
		main_genericstandalone_crc32_checker_syncfifo_consume <= 3'd0;
		main_genericstandalone_rx_converter_converter_source_eop <= 1'd0;
		main_genericstandalone_rx_converter_converter_source_payload_data <= 40'd0;
		main_genericstandalone_rx_converter_converter_demux <= 2'd0;
		main_genericstandalone_rx_converter_converter_strobe_all <= 1'd0;
		main_genericstandalone_rx_cdc_graycounter0_q <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter0_q_binary <= 7'd0;
		builder_a7_1000basex_receivepath_state <= 3'd0;
		builder_liteethmacpreamblechecker_state <= 1'd0;
		builder_liteethmaccrc32checker_state <= 2'd0;
	end
	builder_xilinxmultiregimpl12_regs0 <= main_genericstandalone_rx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl12_regs1 <= builder_xilinxmultiregimpl12_regs0;
end

always @(posedge eth_rx_half_clk) begin
	main_genericstandalone_phase_half_rereg <= main_genericstandalone_phase_half;
end

always @(posedge eth_tx_clk) begin
	main_genericstandalone_pcs_checker_tick <= 1'd0;
	if ((main_genericstandalone_pcs_checker_counter == 1'd0)) begin
		main_genericstandalone_pcs_checker_tick <= 1'd1;
		main_genericstandalone_pcs_checker_counter <= 20'd750000;
	end else begin
		main_genericstandalone_pcs_checker_counter <= (main_genericstandalone_pcs_checker_counter - 1'd1);
	end
	if (main_genericstandalone_pcs_seen_valid_ci_o) begin
		main_genericstandalone_pcs_checker_ok <= 1'd1;
	end
	if (main_genericstandalone_pcs_checker_tick) begin
		main_genericstandalone_pcs_checker_ok <= 1'd0;
	end
	main_genericstandalone_pcs_transmitpath_parity <= (~main_genericstandalone_pcs_transmitpath_parity);
	if (main_genericstandalone_pcs_transmitpath_load_config_reg_buffer) begin
		main_genericstandalone_pcs_transmitpath_config_reg_buffer <= main_genericstandalone_pcs_transmitpath_config_reg;
	end
	main_genericstandalone_pcs_transmitpath_disp_in <= main_genericstandalone_pcs_transmitpath_disp_out;
	main_genericstandalone_pcs_transmitpath_output0 <= main_genericstandalone_pcs_transmitpath_output1;
	main_genericstandalone_pcs_transmitpath_disparity <= main_genericstandalone_pcs_transmitpath_disp_out;
	if ((main_genericstandalone_pcs_transmitpath_k1 & (main_genericstandalone_pcs_transmitpath_d1[4:0] == 5'd28))) begin
		main_genericstandalone_pcs_transmitpath_code6b <= 6'd48;
		main_genericstandalone_pcs_transmitpath_code6b_unbalanced <= 1'd1;
		main_genericstandalone_pcs_transmitpath_code6b_flip <= 1'd1;
	end else begin
		main_genericstandalone_pcs_transmitpath_code6b <= builder_sync_f_rhs_array_muxed1;
		main_genericstandalone_pcs_transmitpath_code6b_unbalanced <= builder_sync_f_rhs_array_muxed2;
		main_genericstandalone_pcs_transmitpath_code6b_flip <= builder_sync_f_rhs_array_muxed3;
	end
	main_genericstandalone_pcs_transmitpath_code4b <= builder_sync_rhs_array_muxed1;
	main_genericstandalone_pcs_transmitpath_code4b_unbalanced <= builder_sync_rhs_array_muxed2;
	if (main_genericstandalone_pcs_transmitpath_k1) begin
		main_genericstandalone_pcs_transmitpath_code4b_flip <= 1'd1;
	end else begin
		main_genericstandalone_pcs_transmitpath_code4b_flip <= builder_sync_f_rhs_array_muxed4;
	end
	main_genericstandalone_pcs_transmitpath_alt7_rd0 <= 1'd0;
	main_genericstandalone_pcs_transmitpath_alt7_rd1 <= 1'd0;
	if ((main_genericstandalone_pcs_transmitpath_d1[7:5] == 3'd7)) begin
		if ((((main_genericstandalone_pcs_transmitpath_d1[4:0] == 5'd17) | (main_genericstandalone_pcs_transmitpath_d1[4:0] == 5'd18)) | (main_genericstandalone_pcs_transmitpath_d1[4:0] == 5'd20))) begin
			main_genericstandalone_pcs_transmitpath_alt7_rd0 <= 1'd1;
		end
		if ((((main_genericstandalone_pcs_transmitpath_d1[4:0] == 4'd11) | (main_genericstandalone_pcs_transmitpath_d1[4:0] == 4'd13)) | (main_genericstandalone_pcs_transmitpath_d1[4:0] == 4'd14))) begin
			main_genericstandalone_pcs_transmitpath_alt7_rd1 <= 1'd1;
		end
		if (main_genericstandalone_pcs_transmitpath_k1) begin
			main_genericstandalone_pcs_transmitpath_alt7_rd0 <= 1'd1;
			main_genericstandalone_pcs_transmitpath_alt7_rd1 <= 1'd1;
		end
	end
	builder_a7_1000basex_transmitpath_state <= builder_a7_1000basex_transmitpath_next_state;
	if (main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value_ce) begin
		main_genericstandalone_pcs_transmitpath_c_type <= main_genericstandalone_pcs_transmitpath_c_type_pcs_next_value;
	end
	main_genericstandalone_pcs_seen_valid_ci_toggle_o_r <= main_genericstandalone_pcs_seen_valid_ci_toggle_o;
	main_genericstandalone_pcs_rx_config_reg_toggle_o_r <= main_genericstandalone_pcs_rx_config_reg_toggle_o;
	main_genericstandalone_pcs_rx_config_reg_ack_toggle_o_r <= main_genericstandalone_pcs_rx_config_reg_ack_toggle_o;
	if (main_genericstandalone_pcs_wait) begin
		if ((~main_genericstandalone_pcs_done)) begin
			main_genericstandalone_pcs_count <= (main_genericstandalone_pcs_count - 1'd1);
		end
	end else begin
		main_genericstandalone_pcs_count <= 21'd1250000;
	end
	builder_a7_1000basex_fsm_state <= builder_a7_1000basex_fsm_next_state;
	if (main_genericstandalone_i) begin
		main_genericstandalone_toggle_i <= (~main_genericstandalone_toggle_i);
	end
	main_genericstandalone_buf <= {main_genericstandalone_tx_data1, main_genericstandalone_buf[19:10]};
	if (main_genericstandalone_tx_gap_inserter_counter_reset) begin
		main_genericstandalone_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_tx_gap_inserter_counter_ce) begin
			main_genericstandalone_tx_gap_inserter_counter <= (main_genericstandalone_tx_gap_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacgap_state <= builder_liteethmacgap_next_state;
	if (main_genericstandalone_preamble_inserter_clr_cnt) begin
		main_genericstandalone_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (main_genericstandalone_preamble_inserter_inc_cnt) begin
			main_genericstandalone_preamble_inserter_cnt <= (main_genericstandalone_preamble_inserter_cnt + 1'd1);
		end
	end
	builder_liteethmacpreambleinserter_state <= builder_liteethmacpreambleinserter_next_state;
	if (main_genericstandalone_crc32_inserter_is_ongoing0) begin
		main_genericstandalone_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((main_genericstandalone_crc32_inserter_is_ongoing1 & (~main_genericstandalone_crc32_inserter_cnt_done))) begin
			main_genericstandalone_crc32_inserter_cnt <= (main_genericstandalone_crc32_inserter_cnt - main_genericstandalone_crc32_inserter_source_ack);
		end
	end
	if (main_genericstandalone_crc32_inserter_ce) begin
		main_genericstandalone_crc32_inserter_reg <= main_genericstandalone_crc32_inserter_next;
	end
	if (main_genericstandalone_crc32_inserter_reset) begin
		main_genericstandalone_crc32_inserter_reg <= 32'd4294967295;
	end
	builder_liteethmaccrc32inserter_state <= builder_liteethmaccrc32inserter_next_state;
	if (main_genericstandalone_padding_inserter_counter_reset) begin
		main_genericstandalone_padding_inserter_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_padding_inserter_counter_ce) begin
			main_genericstandalone_padding_inserter_counter <= (main_genericstandalone_padding_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacpaddinginserter_state <= builder_liteethmacpaddinginserter_next_state;
	if ((main_genericstandalone_tx_last_be_sink_stb & main_genericstandalone_tx_last_be_sink_ack)) begin
		if (main_genericstandalone_tx_last_be_sink_eop) begin
			main_genericstandalone_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (main_genericstandalone_tx_last_be_sink_payload_last_be) begin
				main_genericstandalone_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((main_genericstandalone_tx_converter_converter_source_stb & main_genericstandalone_tx_converter_converter_source_ack)) begin
		if (main_genericstandalone_tx_converter_converter_last) begin
			main_genericstandalone_tx_converter_converter_mux <= 1'd0;
		end else begin
			main_genericstandalone_tx_converter_converter_mux <= (main_genericstandalone_tx_converter_converter_mux + 1'd1);
		end
	end
	main_genericstandalone_tx_cdc_graycounter1_q_binary <= main_genericstandalone_tx_cdc_graycounter1_q_next_binary;
	main_genericstandalone_tx_cdc_graycounter1_q <= main_genericstandalone_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		main_genericstandalone_pcs_transmitpath_output0 <= 10'd0;
		main_genericstandalone_pcs_transmitpath_disparity <= 1'd0;
		main_genericstandalone_pcs_transmitpath_disp_in <= 1'd0;
		main_genericstandalone_pcs_transmitpath_code6b <= 6'd0;
		main_genericstandalone_pcs_transmitpath_code6b_unbalanced <= 1'd0;
		main_genericstandalone_pcs_transmitpath_code6b_flip <= 1'd0;
		main_genericstandalone_pcs_transmitpath_code4b <= 4'd0;
		main_genericstandalone_pcs_transmitpath_code4b_unbalanced <= 1'd0;
		main_genericstandalone_pcs_transmitpath_code4b_flip <= 1'd0;
		main_genericstandalone_pcs_transmitpath_alt7_rd0 <= 1'd0;
		main_genericstandalone_pcs_transmitpath_alt7_rd1 <= 1'd0;
		main_genericstandalone_pcs_transmitpath_parity <= 1'd0;
		main_genericstandalone_pcs_transmitpath_c_type <= 1'd0;
		main_genericstandalone_pcs_transmitpath_config_reg_buffer <= 16'd0;
		main_genericstandalone_pcs_checker_counter <= 20'd0;
		main_genericstandalone_pcs_checker_tick <= 1'd0;
		main_genericstandalone_pcs_checker_ok <= 1'd0;
		main_genericstandalone_pcs_count <= 21'd1250000;
		main_genericstandalone_buf <= 20'd0;
		main_genericstandalone_tx_gap_inserter_counter <= 4'd0;
		main_genericstandalone_preamble_inserter_cnt <= 3'd0;
		main_genericstandalone_crc32_inserter_reg <= 32'd4294967295;
		main_genericstandalone_crc32_inserter_cnt <= 2'd3;
		main_genericstandalone_padding_inserter_counter <= 16'd1;
		main_genericstandalone_tx_last_be_ongoing <= 1'd1;
		main_genericstandalone_tx_converter_converter_mux <= 2'd0;
		main_genericstandalone_tx_cdc_graycounter1_q <= 7'd0;
		main_genericstandalone_tx_cdc_graycounter1_q_binary <= 7'd0;
		builder_a7_1000basex_transmitpath_state <= 3'd0;
		builder_a7_1000basex_fsm_state <= 2'd0;
		builder_liteethmacgap_state <= 1'd0;
		builder_liteethmacpreambleinserter_state <= 2'd0;
		builder_liteethmaccrc32inserter_state <= 2'd0;
		builder_liteethmacpaddinginserter_state <= 1'd0;
	end
	builder_xilinxmultiregimpl1_regs0 <= main_genericstandalone_pcs_seen_valid_ci_toggle_i;
	builder_xilinxmultiregimpl1_regs1 <= builder_xilinxmultiregimpl1_regs0;
	builder_xilinxmultiregimpl2_regs0 <= main_genericstandalone_pcs_rx_config_reg_toggle_i;
	builder_xilinxmultiregimpl2_regs1 <= builder_xilinxmultiregimpl2_regs0;
	builder_xilinxmultiregimpl3_regs0 <= main_genericstandalone_pcs_rx_config_reg_ack_toggle_i;
	builder_xilinxmultiregimpl3_regs1 <= builder_xilinxmultiregimpl3_regs0;
	builder_xilinxmultiregimpl9_regs0 <= main_genericstandalone_tx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl9_regs1 <= builder_xilinxmultiregimpl9_regs0;
end

always @(posedge eth_tx_half_clk) begin
	main_genericstandalone_tx_data_half <= main_genericstandalone_buf;
end

always @(posedge rio_clk) begin
	main_inout_8x0_inout_8x0_sample <= 1'd0;
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & main_inout_8x0_inout_8x0_ointerface0_address[1])) begin
		main_inout_8x0_inout_8x0_sensitivity <= main_inout_8x0_inout_8x0_ointerface0_data;
		if (main_inout_8x0_inout_8x0_ointerface0_address[0]) begin
			main_inout_8x0_inout_8x0_sample <= 1'd1;
		end
	end
	main_inout_8x1_inout_8x1_sample <= 1'd0;
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & main_inout_8x1_inout_8x1_ointerface1_address[1])) begin
		main_inout_8x1_inout_8x1_sensitivity <= main_inout_8x1_inout_8x1_ointerface1_data;
		if (main_inout_8x1_inout_8x1_ointerface1_address[0]) begin
			main_inout_8x1_inout_8x1_sample <= 1'd1;
		end
	end
	main_inout_8x2_inout_8x2_sample <= 1'd0;
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & main_inout_8x2_inout_8x2_ointerface2_address[1])) begin
		main_inout_8x2_inout_8x2_sensitivity <= main_inout_8x2_inout_8x2_ointerface2_data;
		if (main_inout_8x2_inout_8x2_ointerface2_address[0]) begin
			main_inout_8x2_inout_8x2_sample <= 1'd1;
		end
	end
	main_inout_8x3_inout_8x3_sample <= 1'd0;
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & main_inout_8x3_inout_8x3_ointerface3_address[1])) begin
		main_inout_8x3_inout_8x3_sensitivity <= main_inout_8x3_inout_8x3_ointerface3_data;
		if (main_inout_8x3_inout_8x3_ointerface3_address[0]) begin
			main_inout_8x3_inout_8x3_sample <= 1'd1;
		end
	end
	main_inout_8x4_inout_8x4_sample <= 1'd0;
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & main_inout_8x4_inout_8x4_ointerface4_address[1])) begin
		main_inout_8x4_inout_8x4_sensitivity <= main_inout_8x4_inout_8x4_ointerface4_data;
		if (main_inout_8x4_inout_8x4_ointerface4_address[0]) begin
			main_inout_8x4_inout_8x4_sample <= 1'd1;
		end
	end
	main_inout_8x5_inout_8x5_sample <= 1'd0;
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & main_inout_8x5_inout_8x5_ointerface5_address[1])) begin
		main_inout_8x5_inout_8x5_sensitivity <= main_inout_8x5_inout_8x5_ointerface5_data;
		if (main_inout_8x5_inout_8x5_ointerface5_address[0]) begin
			main_inout_8x5_inout_8x5_sample <= 1'd1;
		end
	end
	main_inout_8x6_inout_8x6_sample <= 1'd0;
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & main_inout_8x6_inout_8x6_ointerface6_address[1])) begin
		main_inout_8x6_inout_8x6_sensitivity <= main_inout_8x6_inout_8x6_ointerface6_data;
		if (main_inout_8x6_inout_8x6_ointerface6_address[0]) begin
			main_inout_8x6_inout_8x6_sample <= 1'd1;
		end
	end
	main_inout_8x7_inout_8x7_sample <= 1'd0;
	if ((main_inout_8x7_inout_8x7_ointerface7_stb & main_inout_8x7_inout_8x7_ointerface7_address[1])) begin
		main_inout_8x7_inout_8x7_sensitivity <= main_inout_8x7_inout_8x7_ointerface7_data;
		if (main_inout_8x7_inout_8x7_ointerface7_address[0]) begin
			main_inout_8x7_inout_8x7_sample <= 1'd1;
		end
	end
	if ((main_rtio_core_outputs_asyncfifobuffered0_re | (~main_rtio_core_outputs_asyncfifobuffered0_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered0_dout <= main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
		main_rtio_core_outputs_asyncfifobuffered0_readable <= main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered1_re | (~main_rtio_core_outputs_asyncfifobuffered1_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered1_dout <= main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
		main_rtio_core_outputs_asyncfifobuffered1_readable <= main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered2_re | (~main_rtio_core_outputs_asyncfifobuffered2_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered2_dout <= main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
		main_rtio_core_outputs_asyncfifobuffered2_readable <= main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered3_re | (~main_rtio_core_outputs_asyncfifobuffered3_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered3_dout <= main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
		main_rtio_core_outputs_asyncfifobuffered3_readable <= main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered4_re | (~main_rtio_core_outputs_asyncfifobuffered4_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered4_dout <= main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
		main_rtio_core_outputs_asyncfifobuffered4_readable <= main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered5_re | (~main_rtio_core_outputs_asyncfifobuffered5_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered5_dout <= main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
		main_rtio_core_outputs_asyncfifobuffered5_readable <= main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered6_re | (~main_rtio_core_outputs_asyncfifobuffered6_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered6_dout <= main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
		main_rtio_core_outputs_asyncfifobuffered6_readable <= main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered7_re | (~main_rtio_core_outputs_asyncfifobuffered7_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered7_dout <= main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
		main_rtio_core_outputs_asyncfifobuffered7_readable <= main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
	main_rtio_core_outputs_gates_record0_payload_channel1 <= main_rtio_core_outputs_gates_record0_payload_channel0;
	main_rtio_core_outputs_gates_record0_payload_fine_ts <= main_rtio_core_outputs_gates_record0_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record0_payload_address1 <= main_rtio_core_outputs_gates_record0_payload_address0;
	main_rtio_core_outputs_gates_record0_payload_data1 <= main_rtio_core_outputs_gates_record0_payload_data0;
	main_rtio_core_outputs_gates_record0_seqn1 <= main_rtio_core_outputs_gates_record0_seqn0;
	main_rtio_core_outputs_gates_record0_valid <= (main_rtio_core_outputs_gates_record0_re & main_rtio_core_outputs_gates_record0_readable);
	main_rtio_core_outputs_gates_record1_payload_channel1 <= main_rtio_core_outputs_gates_record1_payload_channel0;
	main_rtio_core_outputs_gates_record1_payload_fine_ts <= main_rtio_core_outputs_gates_record1_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record1_payload_address1 <= main_rtio_core_outputs_gates_record1_payload_address0;
	main_rtio_core_outputs_gates_record1_payload_data1 <= main_rtio_core_outputs_gates_record1_payload_data0;
	main_rtio_core_outputs_gates_record1_seqn1 <= main_rtio_core_outputs_gates_record1_seqn0;
	main_rtio_core_outputs_gates_record1_valid <= (main_rtio_core_outputs_gates_record1_re & main_rtio_core_outputs_gates_record1_readable);
	main_rtio_core_outputs_gates_record2_payload_channel1 <= main_rtio_core_outputs_gates_record2_payload_channel0;
	main_rtio_core_outputs_gates_record2_payload_fine_ts <= main_rtio_core_outputs_gates_record2_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record2_payload_address1 <= main_rtio_core_outputs_gates_record2_payload_address0;
	main_rtio_core_outputs_gates_record2_payload_data1 <= main_rtio_core_outputs_gates_record2_payload_data0;
	main_rtio_core_outputs_gates_record2_seqn1 <= main_rtio_core_outputs_gates_record2_seqn0;
	main_rtio_core_outputs_gates_record2_valid <= (main_rtio_core_outputs_gates_record2_re & main_rtio_core_outputs_gates_record2_readable);
	main_rtio_core_outputs_gates_record3_payload_channel1 <= main_rtio_core_outputs_gates_record3_payload_channel0;
	main_rtio_core_outputs_gates_record3_payload_fine_ts <= main_rtio_core_outputs_gates_record3_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record3_payload_address1 <= main_rtio_core_outputs_gates_record3_payload_address0;
	main_rtio_core_outputs_gates_record3_payload_data1 <= main_rtio_core_outputs_gates_record3_payload_data0;
	main_rtio_core_outputs_gates_record3_seqn1 <= main_rtio_core_outputs_gates_record3_seqn0;
	main_rtio_core_outputs_gates_record3_valid <= (main_rtio_core_outputs_gates_record3_re & main_rtio_core_outputs_gates_record3_readable);
	main_rtio_core_outputs_gates_record4_payload_channel1 <= main_rtio_core_outputs_gates_record4_payload_channel0;
	main_rtio_core_outputs_gates_record4_payload_fine_ts <= main_rtio_core_outputs_gates_record4_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record4_payload_address1 <= main_rtio_core_outputs_gates_record4_payload_address0;
	main_rtio_core_outputs_gates_record4_payload_data1 <= main_rtio_core_outputs_gates_record4_payload_data0;
	main_rtio_core_outputs_gates_record4_seqn1 <= main_rtio_core_outputs_gates_record4_seqn0;
	main_rtio_core_outputs_gates_record4_valid <= (main_rtio_core_outputs_gates_record4_re & main_rtio_core_outputs_gates_record4_readable);
	main_rtio_core_outputs_gates_record5_payload_channel1 <= main_rtio_core_outputs_gates_record5_payload_channel0;
	main_rtio_core_outputs_gates_record5_payload_fine_ts <= main_rtio_core_outputs_gates_record5_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record5_payload_address1 <= main_rtio_core_outputs_gates_record5_payload_address0;
	main_rtio_core_outputs_gates_record5_payload_data1 <= main_rtio_core_outputs_gates_record5_payload_data0;
	main_rtio_core_outputs_gates_record5_seqn1 <= main_rtio_core_outputs_gates_record5_seqn0;
	main_rtio_core_outputs_gates_record5_valid <= (main_rtio_core_outputs_gates_record5_re & main_rtio_core_outputs_gates_record5_readable);
	main_rtio_core_outputs_gates_record6_payload_channel1 <= main_rtio_core_outputs_gates_record6_payload_channel0;
	main_rtio_core_outputs_gates_record6_payload_fine_ts <= main_rtio_core_outputs_gates_record6_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record6_payload_address1 <= main_rtio_core_outputs_gates_record6_payload_address0;
	main_rtio_core_outputs_gates_record6_payload_data1 <= main_rtio_core_outputs_gates_record6_payload_data0;
	main_rtio_core_outputs_gates_record6_seqn1 <= main_rtio_core_outputs_gates_record6_seqn0;
	main_rtio_core_outputs_gates_record6_valid <= (main_rtio_core_outputs_gates_record6_re & main_rtio_core_outputs_gates_record6_readable);
	main_rtio_core_outputs_gates_record7_payload_channel1 <= main_rtio_core_outputs_gates_record7_payload_channel0;
	main_rtio_core_outputs_gates_record7_payload_fine_ts <= main_rtio_core_outputs_gates_record7_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record7_payload_address1 <= main_rtio_core_outputs_gates_record7_payload_address0;
	main_rtio_core_outputs_gates_record7_payload_data1 <= main_rtio_core_outputs_gates_record7_payload_data0;
	main_rtio_core_outputs_gates_record7_seqn1 <= main_rtio_core_outputs_gates_record7_seqn0;
	main_rtio_core_outputs_gates_record7_valid <= (main_rtio_core_outputs_gates_record7_re & main_rtio_core_outputs_gates_record7_readable);
	main_rtio_core_outputs_record0_valid1 <= main_rtio_core_outputs_record40_rec_valid;
	main_rtio_core_outputs_record0_payload_channel3 <= main_rtio_core_outputs_record40_rec_payload_channel;
	main_rtio_core_outputs_record0_payload_fine_ts1 <= main_rtio_core_outputs_record40_rec_payload_fine_ts;
	main_rtio_core_outputs_record0_payload_address3 <= main_rtio_core_outputs_record40_rec_payload_address;
	main_rtio_core_outputs_record0_payload_data3 <= main_rtio_core_outputs_record40_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r0 <= main_rtio_core_outputs_record40_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r0 <= main_rtio_core_outputs_record40_rec_nondata_replace_occured;
	main_rtio_core_outputs_record1_valid1 <= main_rtio_core_outputs_record41_rec_valid;
	main_rtio_core_outputs_record1_payload_channel3 <= main_rtio_core_outputs_record41_rec_payload_channel;
	main_rtio_core_outputs_record1_payload_fine_ts1 <= main_rtio_core_outputs_record41_rec_payload_fine_ts;
	main_rtio_core_outputs_record1_payload_address3 <= main_rtio_core_outputs_record41_rec_payload_address;
	main_rtio_core_outputs_record1_payload_data3 <= main_rtio_core_outputs_record41_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r1 <= main_rtio_core_outputs_record41_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r1 <= main_rtio_core_outputs_record41_rec_nondata_replace_occured;
	main_rtio_core_outputs_record2_valid1 <= main_rtio_core_outputs_record42_rec_valid;
	main_rtio_core_outputs_record2_payload_channel3 <= main_rtio_core_outputs_record42_rec_payload_channel;
	main_rtio_core_outputs_record2_payload_fine_ts1 <= main_rtio_core_outputs_record42_rec_payload_fine_ts;
	main_rtio_core_outputs_record2_payload_address3 <= main_rtio_core_outputs_record42_rec_payload_address;
	main_rtio_core_outputs_record2_payload_data3 <= main_rtio_core_outputs_record42_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r2 <= main_rtio_core_outputs_record42_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r2 <= main_rtio_core_outputs_record42_rec_nondata_replace_occured;
	main_rtio_core_outputs_record3_valid1 <= main_rtio_core_outputs_record43_rec_valid;
	main_rtio_core_outputs_record3_payload_channel3 <= main_rtio_core_outputs_record43_rec_payload_channel;
	main_rtio_core_outputs_record3_payload_fine_ts1 <= main_rtio_core_outputs_record43_rec_payload_fine_ts;
	main_rtio_core_outputs_record3_payload_address3 <= main_rtio_core_outputs_record43_rec_payload_address;
	main_rtio_core_outputs_record3_payload_data3 <= main_rtio_core_outputs_record43_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r3 <= main_rtio_core_outputs_record43_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r3 <= main_rtio_core_outputs_record43_rec_nondata_replace_occured;
	main_rtio_core_outputs_record4_valid1 <= main_rtio_core_outputs_record44_rec_valid;
	main_rtio_core_outputs_record4_payload_channel3 <= main_rtio_core_outputs_record44_rec_payload_channel;
	main_rtio_core_outputs_record4_payload_fine_ts1 <= main_rtio_core_outputs_record44_rec_payload_fine_ts;
	main_rtio_core_outputs_record4_payload_address3 <= main_rtio_core_outputs_record44_rec_payload_address;
	main_rtio_core_outputs_record4_payload_data3 <= main_rtio_core_outputs_record44_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r4 <= main_rtio_core_outputs_record44_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r4 <= main_rtio_core_outputs_record44_rec_nondata_replace_occured;
	main_rtio_core_outputs_record5_valid1 <= main_rtio_core_outputs_record45_rec_valid;
	main_rtio_core_outputs_record5_payload_channel3 <= main_rtio_core_outputs_record45_rec_payload_channel;
	main_rtio_core_outputs_record5_payload_fine_ts1 <= main_rtio_core_outputs_record45_rec_payload_fine_ts;
	main_rtio_core_outputs_record5_payload_address3 <= main_rtio_core_outputs_record45_rec_payload_address;
	main_rtio_core_outputs_record5_payload_data3 <= main_rtio_core_outputs_record45_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r5 <= main_rtio_core_outputs_record45_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r5 <= main_rtio_core_outputs_record45_rec_nondata_replace_occured;
	main_rtio_core_outputs_record6_valid1 <= main_rtio_core_outputs_record46_rec_valid;
	main_rtio_core_outputs_record6_payload_channel3 <= main_rtio_core_outputs_record46_rec_payload_channel;
	main_rtio_core_outputs_record6_payload_fine_ts1 <= main_rtio_core_outputs_record46_rec_payload_fine_ts;
	main_rtio_core_outputs_record6_payload_address3 <= main_rtio_core_outputs_record46_rec_payload_address;
	main_rtio_core_outputs_record6_payload_data3 <= main_rtio_core_outputs_record46_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r6 <= main_rtio_core_outputs_record46_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r6 <= main_rtio_core_outputs_record46_rec_nondata_replace_occured;
	main_rtio_core_outputs_record7_valid1 <= main_rtio_core_outputs_record47_rec_valid;
	main_rtio_core_outputs_record7_payload_channel3 <= main_rtio_core_outputs_record47_rec_payload_channel;
	main_rtio_core_outputs_record7_payload_fine_ts1 <= main_rtio_core_outputs_record47_rec_payload_fine_ts;
	main_rtio_core_outputs_record7_payload_address3 <= main_rtio_core_outputs_record47_rec_payload_address;
	main_rtio_core_outputs_record7_payload_data3 <= main_rtio_core_outputs_record47_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r7 <= main_rtio_core_outputs_record47_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r7 <= main_rtio_core_outputs_record47_rec_nondata_replace_occured;
	main_rtio_core_outputs_collision <= 1'd0;
	main_rtio_core_outputs_collision_channel <= 1'd0;
	if ((main_rtio_core_outputs_record0_valid1 & main_rtio_core_outputs_record0_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record0_payload_channel3;
	end
	if ((main_rtio_core_outputs_record1_valid1 & main_rtio_core_outputs_record1_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record1_payload_channel3;
	end
	if ((main_rtio_core_outputs_record2_valid1 & main_rtio_core_outputs_record2_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record2_payload_channel3;
	end
	if ((main_rtio_core_outputs_record3_valid1 & main_rtio_core_outputs_record3_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record3_payload_channel3;
	end
	if ((main_rtio_core_outputs_record4_valid1 & main_rtio_core_outputs_record4_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record4_payload_channel3;
	end
	if ((main_rtio_core_outputs_record5_valid1 & main_rtio_core_outputs_record5_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record5_payload_channel3;
	end
	if ((main_rtio_core_outputs_record6_valid1 & main_rtio_core_outputs_record6_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record6_payload_channel3;
	end
	if ((main_rtio_core_outputs_record7_valid1 & main_rtio_core_outputs_record7_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record7_payload_channel3;
	end
	main_inout_8x0_inout_8x0_ointerface0_stb <= (((((((main_rtio_core_outputs_selected0 | main_rtio_core_outputs_selected1) | main_rtio_core_outputs_selected2) | main_rtio_core_outputs_selected3) | main_rtio_core_outputs_selected4) | main_rtio_core_outputs_selected5) | main_rtio_core_outputs_selected6) | main_rtio_core_outputs_selected7);
	main_inout_8x0_inout_8x0_ointerface0_fine_ts <= ((((((((main_rtio_core_outputs_selected0 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected1 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected2 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected3 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected4 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected5 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected6 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected7 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_address <= ((((((((main_rtio_core_outputs_selected0 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected1 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected2 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected3 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected4 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected5 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected6 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected7 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_data <= ((((((((main_rtio_core_outputs_selected0 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected1 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected2 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected3 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected4 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected5 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected6 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected7 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_stb <= (((((((main_rtio_core_outputs_selected8 | main_rtio_core_outputs_selected9) | main_rtio_core_outputs_selected10) | main_rtio_core_outputs_selected11) | main_rtio_core_outputs_selected12) | main_rtio_core_outputs_selected13) | main_rtio_core_outputs_selected14) | main_rtio_core_outputs_selected15);
	main_inout_8x1_inout_8x1_ointerface1_fine_ts <= ((((((((main_rtio_core_outputs_selected8 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected9 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected10 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected11 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected12 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected13 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected14 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected15 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_address <= ((((((((main_rtio_core_outputs_selected8 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected9 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected10 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected11 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected12 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected13 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected14 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected15 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_data <= ((((((((main_rtio_core_outputs_selected8 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected9 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected10 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected11 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected12 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected13 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected14 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected15 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_stb <= (((((((main_rtio_core_outputs_selected16 | main_rtio_core_outputs_selected17) | main_rtio_core_outputs_selected18) | main_rtio_core_outputs_selected19) | main_rtio_core_outputs_selected20) | main_rtio_core_outputs_selected21) | main_rtio_core_outputs_selected22) | main_rtio_core_outputs_selected23);
	main_inout_8x2_inout_8x2_ointerface2_fine_ts <= ((((((((main_rtio_core_outputs_selected16 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected17 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected18 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected19 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected20 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected21 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected22 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected23 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_address <= ((((((((main_rtio_core_outputs_selected16 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected17 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected18 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected19 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected20 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected21 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected22 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected23 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_data <= ((((((((main_rtio_core_outputs_selected16 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected17 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected18 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected19 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected20 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected21 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected22 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected23 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_stb <= (((((((main_rtio_core_outputs_selected24 | main_rtio_core_outputs_selected25) | main_rtio_core_outputs_selected26) | main_rtio_core_outputs_selected27) | main_rtio_core_outputs_selected28) | main_rtio_core_outputs_selected29) | main_rtio_core_outputs_selected30) | main_rtio_core_outputs_selected31);
	main_inout_8x3_inout_8x3_ointerface3_fine_ts <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_address <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_data <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_stb <= (((((((main_rtio_core_outputs_selected32 | main_rtio_core_outputs_selected33) | main_rtio_core_outputs_selected34) | main_rtio_core_outputs_selected35) | main_rtio_core_outputs_selected36) | main_rtio_core_outputs_selected37) | main_rtio_core_outputs_selected38) | main_rtio_core_outputs_selected39);
	main_inout_8x4_inout_8x4_ointerface4_fine_ts <= ((((((((main_rtio_core_outputs_selected32 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected33 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected34 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected35 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected36 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected37 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected38 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected39 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_address <= ((((((((main_rtio_core_outputs_selected32 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected33 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected34 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected35 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected36 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected37 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected38 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected39 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_data <= ((((((((main_rtio_core_outputs_selected32 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected33 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected34 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected35 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected36 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected37 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected38 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected39 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_stb <= (((((((main_rtio_core_outputs_selected40 | main_rtio_core_outputs_selected41) | main_rtio_core_outputs_selected42) | main_rtio_core_outputs_selected43) | main_rtio_core_outputs_selected44) | main_rtio_core_outputs_selected45) | main_rtio_core_outputs_selected46) | main_rtio_core_outputs_selected47);
	main_inout_8x5_inout_8x5_ointerface5_fine_ts <= ((((((((main_rtio_core_outputs_selected40 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected41 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected42 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected43 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected44 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected45 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected46 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected47 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_address <= ((((((((main_rtio_core_outputs_selected40 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected41 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected42 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected43 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected44 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected45 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected46 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected47 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_data <= ((((((((main_rtio_core_outputs_selected40 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected41 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected42 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected43 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected44 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected45 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected46 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected47 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_stb <= (((((((main_rtio_core_outputs_selected48 | main_rtio_core_outputs_selected49) | main_rtio_core_outputs_selected50) | main_rtio_core_outputs_selected51) | main_rtio_core_outputs_selected52) | main_rtio_core_outputs_selected53) | main_rtio_core_outputs_selected54) | main_rtio_core_outputs_selected55);
	main_inout_8x6_inout_8x6_ointerface6_fine_ts <= ((((((((main_rtio_core_outputs_selected48 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected49 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected50 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected51 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected52 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected53 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected54 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected55 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_address <= ((((((((main_rtio_core_outputs_selected48 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected49 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected50 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected51 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected52 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected53 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected54 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected55 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_data <= ((((((((main_rtio_core_outputs_selected48 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected49 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected50 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected51 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected52 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected53 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected54 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected55 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x7_inout_8x7_ointerface7_stb <= (((((((main_rtio_core_outputs_selected56 | main_rtio_core_outputs_selected57) | main_rtio_core_outputs_selected58) | main_rtio_core_outputs_selected59) | main_rtio_core_outputs_selected60) | main_rtio_core_outputs_selected61) | main_rtio_core_outputs_selected62) | main_rtio_core_outputs_selected63);
	main_inout_8x7_inout_8x7_ointerface7_fine_ts <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x7_inout_8x7_ointerface7_address <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x7_inout_8x7_ointerface7_data <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x0_stb <= (((((((main_rtio_core_outputs_selected64 | main_rtio_core_outputs_selected65) | main_rtio_core_outputs_selected66) | main_rtio_core_outputs_selected67) | main_rtio_core_outputs_selected68) | main_rtio_core_outputs_selected69) | main_rtio_core_outputs_selected70) | main_rtio_core_outputs_selected71);
	main_output_8x0_fine_ts <= ((((((((main_rtio_core_outputs_selected64 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected65 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected66 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected67 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected68 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected69 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected70 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected71 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x0_data <= ((((((((main_rtio_core_outputs_selected64 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected65 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected66 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected67 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected68 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected69 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected70 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected71 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x1_stb <= (((((((main_rtio_core_outputs_selected72 | main_rtio_core_outputs_selected73) | main_rtio_core_outputs_selected74) | main_rtio_core_outputs_selected75) | main_rtio_core_outputs_selected76) | main_rtio_core_outputs_selected77) | main_rtio_core_outputs_selected78) | main_rtio_core_outputs_selected79);
	main_output_8x1_fine_ts <= ((((((((main_rtio_core_outputs_selected72 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected73 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected74 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected75 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected76 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected77 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected78 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected79 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x1_data <= ((((((((main_rtio_core_outputs_selected72 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected73 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected74 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected75 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected76 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected77 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected78 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected79 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x2_stb <= (((((((main_rtio_core_outputs_selected80 | main_rtio_core_outputs_selected81) | main_rtio_core_outputs_selected82) | main_rtio_core_outputs_selected83) | main_rtio_core_outputs_selected84) | main_rtio_core_outputs_selected85) | main_rtio_core_outputs_selected86) | main_rtio_core_outputs_selected87);
	main_output_8x2_fine_ts <= ((((((((main_rtio_core_outputs_selected80 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected81 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected82 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected83 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected84 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected85 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected86 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected87 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x2_data <= ((((((((main_rtio_core_outputs_selected80 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected81 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected82 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected83 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected84 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected85 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected86 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected87 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x3_stb <= (((((((main_rtio_core_outputs_selected88 | main_rtio_core_outputs_selected89) | main_rtio_core_outputs_selected90) | main_rtio_core_outputs_selected91) | main_rtio_core_outputs_selected92) | main_rtio_core_outputs_selected93) | main_rtio_core_outputs_selected94) | main_rtio_core_outputs_selected95);
	main_output_8x3_fine_ts <= ((((((((main_rtio_core_outputs_selected88 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected89 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected90 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected91 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected92 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected93 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected94 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected95 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x3_data <= ((((((((main_rtio_core_outputs_selected88 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected89 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected90 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected91 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected92 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected93 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected94 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected95 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x4_stb <= (((((((main_rtio_core_outputs_selected96 | main_rtio_core_outputs_selected97) | main_rtio_core_outputs_selected98) | main_rtio_core_outputs_selected99) | main_rtio_core_outputs_selected100) | main_rtio_core_outputs_selected101) | main_rtio_core_outputs_selected102) | main_rtio_core_outputs_selected103);
	main_output_8x4_fine_ts <= ((((((((main_rtio_core_outputs_selected96 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected97 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected98 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected99 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected100 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected101 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected102 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected103 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x4_data <= ((((((((main_rtio_core_outputs_selected96 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected97 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected98 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected99 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected100 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected101 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected102 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected103 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x5_stb <= (((((((main_rtio_core_outputs_selected104 | main_rtio_core_outputs_selected105) | main_rtio_core_outputs_selected106) | main_rtio_core_outputs_selected107) | main_rtio_core_outputs_selected108) | main_rtio_core_outputs_selected109) | main_rtio_core_outputs_selected110) | main_rtio_core_outputs_selected111);
	main_output_8x5_fine_ts <= ((((((((main_rtio_core_outputs_selected104 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected105 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected106 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected107 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected108 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected109 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected110 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected111 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x5_data <= ((((((((main_rtio_core_outputs_selected104 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected105 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected106 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected107 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected108 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected109 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected110 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected111 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x6_stb <= (((((((main_rtio_core_outputs_selected112 | main_rtio_core_outputs_selected113) | main_rtio_core_outputs_selected114) | main_rtio_core_outputs_selected115) | main_rtio_core_outputs_selected116) | main_rtio_core_outputs_selected117) | main_rtio_core_outputs_selected118) | main_rtio_core_outputs_selected119);
	main_output_8x6_fine_ts <= ((((((((main_rtio_core_outputs_selected112 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected113 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected114 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected115 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected116 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected117 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected118 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected119 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x6_data <= ((((((((main_rtio_core_outputs_selected112 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected113 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected114 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected115 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected116 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected117 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected118 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected119 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x7_stb <= (((((((main_rtio_core_outputs_selected120 | main_rtio_core_outputs_selected121) | main_rtio_core_outputs_selected122) | main_rtio_core_outputs_selected123) | main_rtio_core_outputs_selected124) | main_rtio_core_outputs_selected125) | main_rtio_core_outputs_selected126) | main_rtio_core_outputs_selected127);
	main_output_8x7_fine_ts <= ((((((((main_rtio_core_outputs_selected120 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected121 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected122 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected123 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected124 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected125 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected126 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected127 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x7_data <= ((((((((main_rtio_core_outputs_selected120 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected121 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected122 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected123 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected124 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected125 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected126 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected127 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster0_ointerface0_stb <= (((((((main_rtio_core_outputs_selected128 | main_rtio_core_outputs_selected129) | main_rtio_core_outputs_selected130) | main_rtio_core_outputs_selected131) | main_rtio_core_outputs_selected132) | main_rtio_core_outputs_selected133) | main_rtio_core_outputs_selected134) | main_rtio_core_outputs_selected135);
	main_spimaster0_ointerface0_address <= ((((((((main_rtio_core_outputs_selected128 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected129 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected130 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected131 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected132 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected133 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected134 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected135 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster0_ointerface0_data <= ((((((((main_rtio_core_outputs_selected128 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected129 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected130 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected131 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected132 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected133 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected134 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected135 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x8_stb <= (((((((main_rtio_core_outputs_selected136 | main_rtio_core_outputs_selected137) | main_rtio_core_outputs_selected138) | main_rtio_core_outputs_selected139) | main_rtio_core_outputs_selected140) | main_rtio_core_outputs_selected141) | main_rtio_core_outputs_selected142) | main_rtio_core_outputs_selected143);
	main_output_8x8_fine_ts <= ((((((((main_rtio_core_outputs_selected136 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected137 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected138 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected139 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected140 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected141 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected142 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected143 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x8_data <= ((((((((main_rtio_core_outputs_selected136 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected137 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected138 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected139 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected140 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected141 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected142 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected143 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x9_stb <= (((((((main_rtio_core_outputs_selected144 | main_rtio_core_outputs_selected145) | main_rtio_core_outputs_selected146) | main_rtio_core_outputs_selected147) | main_rtio_core_outputs_selected148) | main_rtio_core_outputs_selected149) | main_rtio_core_outputs_selected150) | main_rtio_core_outputs_selected151);
	main_output_8x9_fine_ts <= ((((((((main_rtio_core_outputs_selected144 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected145 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected146 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected147 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected148 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected149 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected150 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected151 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x9_data <= ((((((((main_rtio_core_outputs_selected144 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected145 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected146 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected147 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected148 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected149 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected150 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected151 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x10_stb <= (((((((main_rtio_core_outputs_selected152 | main_rtio_core_outputs_selected153) | main_rtio_core_outputs_selected154) | main_rtio_core_outputs_selected155) | main_rtio_core_outputs_selected156) | main_rtio_core_outputs_selected157) | main_rtio_core_outputs_selected158) | main_rtio_core_outputs_selected159);
	main_output_8x10_fine_ts <= ((((((((main_rtio_core_outputs_selected152 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected153 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected154 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected155 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected156 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected157 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected158 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected159 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x10_data <= ((((((((main_rtio_core_outputs_selected152 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected153 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected154 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected155 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected156 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected157 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected158 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected159 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x11_stb <= (((((((main_rtio_core_outputs_selected160 | main_rtio_core_outputs_selected161) | main_rtio_core_outputs_selected162) | main_rtio_core_outputs_selected163) | main_rtio_core_outputs_selected164) | main_rtio_core_outputs_selected165) | main_rtio_core_outputs_selected166) | main_rtio_core_outputs_selected167);
	main_output_8x11_fine_ts <= ((((((((main_rtio_core_outputs_selected160 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected161 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected162 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected163 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected164 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected165 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected166 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected167 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x11_data <= ((((((((main_rtio_core_outputs_selected160 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected161 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected162 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected163 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected164 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected165 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected166 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected167 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x12_stb <= (((((((main_rtio_core_outputs_selected168 | main_rtio_core_outputs_selected169) | main_rtio_core_outputs_selected170) | main_rtio_core_outputs_selected171) | main_rtio_core_outputs_selected172) | main_rtio_core_outputs_selected173) | main_rtio_core_outputs_selected174) | main_rtio_core_outputs_selected175);
	main_output_8x12_fine_ts <= ((((((((main_rtio_core_outputs_selected168 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected169 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected170 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected171 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected172 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected173 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected174 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected175 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x12_data <= ((((((((main_rtio_core_outputs_selected168 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected169 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected170 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected171 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected172 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected173 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected174 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected175 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster1_ointerface1_stb <= (((((((main_rtio_core_outputs_selected176 | main_rtio_core_outputs_selected177) | main_rtio_core_outputs_selected178) | main_rtio_core_outputs_selected179) | main_rtio_core_outputs_selected180) | main_rtio_core_outputs_selected181) | main_rtio_core_outputs_selected182) | main_rtio_core_outputs_selected183);
	main_spimaster1_ointerface1_address <= ((((((((main_rtio_core_outputs_selected176 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected177 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected178 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected179 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected180 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected181 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected182 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected183 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster1_ointerface1_data <= ((((((((main_rtio_core_outputs_selected176 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected177 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected178 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected179 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected180 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected181 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected182 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected183 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x13_stb <= (((((((main_rtio_core_outputs_selected184 | main_rtio_core_outputs_selected185) | main_rtio_core_outputs_selected186) | main_rtio_core_outputs_selected187) | main_rtio_core_outputs_selected188) | main_rtio_core_outputs_selected189) | main_rtio_core_outputs_selected190) | main_rtio_core_outputs_selected191);
	main_output_8x13_fine_ts <= ((((((((main_rtio_core_outputs_selected184 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected185 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected186 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected187 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected188 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected189 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected190 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected191 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x13_data <= ((((((((main_rtio_core_outputs_selected184 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected185 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected186 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected187 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected188 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected189 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected190 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected191 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x14_stb <= (((((((main_rtio_core_outputs_selected192 | main_rtio_core_outputs_selected193) | main_rtio_core_outputs_selected194) | main_rtio_core_outputs_selected195) | main_rtio_core_outputs_selected196) | main_rtio_core_outputs_selected197) | main_rtio_core_outputs_selected198) | main_rtio_core_outputs_selected199);
	main_output_8x14_fine_ts <= ((((((((main_rtio_core_outputs_selected192 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected193 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected194 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected195 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected196 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected197 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected198 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected199 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x14_data <= ((((((((main_rtio_core_outputs_selected192 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected193 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected194 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected195 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected196 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected197 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected198 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected199 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x15_stb <= (((((((main_rtio_core_outputs_selected200 | main_rtio_core_outputs_selected201) | main_rtio_core_outputs_selected202) | main_rtio_core_outputs_selected203) | main_rtio_core_outputs_selected204) | main_rtio_core_outputs_selected205) | main_rtio_core_outputs_selected206) | main_rtio_core_outputs_selected207);
	main_output_8x15_fine_ts <= ((((((((main_rtio_core_outputs_selected200 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected201 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected202 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected203 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected204 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected205 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected206 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected207 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x15_data <= ((((((((main_rtio_core_outputs_selected200 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected201 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected202 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected203 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected204 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected205 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected206 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected207 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x16_stb <= (((((((main_rtio_core_outputs_selected208 | main_rtio_core_outputs_selected209) | main_rtio_core_outputs_selected210) | main_rtio_core_outputs_selected211) | main_rtio_core_outputs_selected212) | main_rtio_core_outputs_selected213) | main_rtio_core_outputs_selected214) | main_rtio_core_outputs_selected215);
	main_output_8x16_fine_ts <= ((((((((main_rtio_core_outputs_selected208 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected209 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected210 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected211 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected212 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected213 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected214 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected215 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x16_data <= ((((((((main_rtio_core_outputs_selected208 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected209 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected210 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected211 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected212 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected213 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected214 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected215 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x17_stb <= (((((((main_rtio_core_outputs_selected216 | main_rtio_core_outputs_selected217) | main_rtio_core_outputs_selected218) | main_rtio_core_outputs_selected219) | main_rtio_core_outputs_selected220) | main_rtio_core_outputs_selected221) | main_rtio_core_outputs_selected222) | main_rtio_core_outputs_selected223);
	main_output_8x17_fine_ts <= ((((((((main_rtio_core_outputs_selected216 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected217 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected218 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected219 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected220 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected221 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected222 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected223 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x17_data <= ((((((((main_rtio_core_outputs_selected216 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected217 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected218 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected219 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected220 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected221 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected222 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected223 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster2_ointerface2_stb <= (((((((main_rtio_core_outputs_selected224 | main_rtio_core_outputs_selected225) | main_rtio_core_outputs_selected226) | main_rtio_core_outputs_selected227) | main_rtio_core_outputs_selected228) | main_rtio_core_outputs_selected229) | main_rtio_core_outputs_selected230) | main_rtio_core_outputs_selected231);
	main_spimaster2_ointerface2_address <= ((((((((main_rtio_core_outputs_selected224 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected225 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected226 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected227 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected228 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected229 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected230 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected231 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster2_ointerface2_data <= ((((((((main_rtio_core_outputs_selected224 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected225 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected226 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected227 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected228 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected229 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected230 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected231 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x18_stb <= (((((((main_rtio_core_outputs_selected232 | main_rtio_core_outputs_selected233) | main_rtio_core_outputs_selected234) | main_rtio_core_outputs_selected235) | main_rtio_core_outputs_selected236) | main_rtio_core_outputs_selected237) | main_rtio_core_outputs_selected238) | main_rtio_core_outputs_selected239);
	main_output_8x18_fine_ts <= ((((((((main_rtio_core_outputs_selected232 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected233 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected234 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected235 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected236 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected237 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected238 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected239 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x18_data <= ((((((((main_rtio_core_outputs_selected232 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected233 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected234 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected235 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected236 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected237 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected238 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected239 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x19_stb <= (((((((main_rtio_core_outputs_selected240 | main_rtio_core_outputs_selected241) | main_rtio_core_outputs_selected242) | main_rtio_core_outputs_selected243) | main_rtio_core_outputs_selected244) | main_rtio_core_outputs_selected245) | main_rtio_core_outputs_selected246) | main_rtio_core_outputs_selected247);
	main_output_8x19_fine_ts <= ((((((((main_rtio_core_outputs_selected240 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected241 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected242 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected243 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected244 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected245 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected246 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected247 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x19_data <= ((((((((main_rtio_core_outputs_selected240 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected241 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected242 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected243 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected244 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected245 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected246 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected247 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x20_stb <= (((((((main_rtio_core_outputs_selected248 | main_rtio_core_outputs_selected249) | main_rtio_core_outputs_selected250) | main_rtio_core_outputs_selected251) | main_rtio_core_outputs_selected252) | main_rtio_core_outputs_selected253) | main_rtio_core_outputs_selected254) | main_rtio_core_outputs_selected255);
	main_output_8x20_fine_ts <= ((((((((main_rtio_core_outputs_selected248 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected249 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected250 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected251 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected252 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected253 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected254 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected255 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x20_data <= ((((((((main_rtio_core_outputs_selected248 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected249 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected250 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected251 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected252 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected253 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected254 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected255 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x21_stb <= (((((((main_rtio_core_outputs_selected256 | main_rtio_core_outputs_selected257) | main_rtio_core_outputs_selected258) | main_rtio_core_outputs_selected259) | main_rtio_core_outputs_selected260) | main_rtio_core_outputs_selected261) | main_rtio_core_outputs_selected262) | main_rtio_core_outputs_selected263);
	main_output_8x21_fine_ts <= ((((((((main_rtio_core_outputs_selected256 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected257 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected258 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected259 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected260 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected261 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected262 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected263 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x21_data <= ((((((((main_rtio_core_outputs_selected256 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected257 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected258 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected259 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected260 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected261 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected262 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected263 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x22_stb <= (((((((main_rtio_core_outputs_selected264 | main_rtio_core_outputs_selected265) | main_rtio_core_outputs_selected266) | main_rtio_core_outputs_selected267) | main_rtio_core_outputs_selected268) | main_rtio_core_outputs_selected269) | main_rtio_core_outputs_selected270) | main_rtio_core_outputs_selected271);
	main_output_8x22_fine_ts <= ((((((((main_rtio_core_outputs_selected264 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected265 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected266 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected267 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected268 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected269 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected270 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected271 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x22_data <= ((((((((main_rtio_core_outputs_selected264 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected265 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected266 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected267 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected268 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected269 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected270 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected271 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output0_stb <= (((((((main_rtio_core_outputs_selected272 | main_rtio_core_outputs_selected273) | main_rtio_core_outputs_selected274) | main_rtio_core_outputs_selected275) | main_rtio_core_outputs_selected276) | main_rtio_core_outputs_selected277) | main_rtio_core_outputs_selected278) | main_rtio_core_outputs_selected279);
	main_output0_data <= ((((((((main_rtio_core_outputs_selected272 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected273 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected274 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected275 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected276 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected277 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected278 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected279 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output1_stb <= (((((((main_rtio_core_outputs_selected280 | main_rtio_core_outputs_selected281) | main_rtio_core_outputs_selected282) | main_rtio_core_outputs_selected283) | main_rtio_core_outputs_selected284) | main_rtio_core_outputs_selected285) | main_rtio_core_outputs_selected286) | main_rtio_core_outputs_selected287);
	main_output1_data <= ((((((((main_rtio_core_outputs_selected280 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected281 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected282 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected283 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected284 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected285 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected286 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected287 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_stb <= (((((((main_rtio_core_outputs_selected288 | main_rtio_core_outputs_selected289) | main_rtio_core_outputs_selected290) | main_rtio_core_outputs_selected291) | main_rtio_core_outputs_selected292) | main_rtio_core_outputs_selected293) | main_rtio_core_outputs_selected294) | main_rtio_core_outputs_selected295);
	main_data <= ((((((((main_rtio_core_outputs_selected288 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected289 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected290 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected291 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected292 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected293 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected294 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected295 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_rtio_core_outputs_busy <= 1'd0;
	main_rtio_core_outputs_busy_channel <= 1'd0;
	main_rtio_core_outputs_stb_r0 <= (main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision));
	main_rtio_core_outputs_channel_r0 <= main_rtio_core_outputs_record0_payload_channel3;
	if ((main_rtio_core_outputs_stb_r0 & builder_sync_basiclowerer_array_muxed0)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r0;
	end
	main_rtio_core_outputs_stb_r1 <= (main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision));
	main_rtio_core_outputs_channel_r1 <= main_rtio_core_outputs_record1_payload_channel3;
	if ((main_rtio_core_outputs_stb_r1 & builder_sync_basiclowerer_array_muxed1)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r1;
	end
	main_rtio_core_outputs_stb_r2 <= (main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision));
	main_rtio_core_outputs_channel_r2 <= main_rtio_core_outputs_record2_payload_channel3;
	if ((main_rtio_core_outputs_stb_r2 & builder_sync_basiclowerer_array_muxed2)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r2;
	end
	main_rtio_core_outputs_stb_r3 <= (main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision));
	main_rtio_core_outputs_channel_r3 <= main_rtio_core_outputs_record3_payload_channel3;
	if ((main_rtio_core_outputs_stb_r3 & builder_sync_basiclowerer_array_muxed3)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r3;
	end
	main_rtio_core_outputs_stb_r4 <= (main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision));
	main_rtio_core_outputs_channel_r4 <= main_rtio_core_outputs_record4_payload_channel3;
	if ((main_rtio_core_outputs_stb_r4 & builder_sync_basiclowerer_array_muxed4)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r4;
	end
	main_rtio_core_outputs_stb_r5 <= (main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision));
	main_rtio_core_outputs_channel_r5 <= main_rtio_core_outputs_record5_payload_channel3;
	if ((main_rtio_core_outputs_stb_r5 & builder_sync_basiclowerer_array_muxed5)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r5;
	end
	main_rtio_core_outputs_stb_r6 <= (main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision));
	main_rtio_core_outputs_channel_r6 <= main_rtio_core_outputs_record6_payload_channel3;
	if ((main_rtio_core_outputs_stb_r6 & builder_sync_basiclowerer_array_muxed6)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r6;
	end
	main_rtio_core_outputs_stb_r7 <= (main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision));
	main_rtio_core_outputs_channel_r7 <= main_rtio_core_outputs_record7_payload_channel3;
	if ((main_rtio_core_outputs_stb_r7 & builder_sync_basiclowerer_array_muxed7)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r7;
	end
	if (({(~main_rtio_core_outputs_record0_valid0), main_rtio_core_outputs_record0_payload_channel2} == {(~main_rtio_core_outputs_record1_valid0), main_rtio_core_outputs_record1_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record0_seqn2[10] == main_rtio_core_outputs_record0_seqn2[11]) & (main_rtio_core_outputs_record1_seqn2[10] == main_rtio_core_outputs_record1_seqn2[11])) & (main_rtio_core_outputs_record0_seqn2[11] != main_rtio_core_outputs_record1_seqn2[11])) ? main_rtio_core_outputs_record0_seqn2[11] : (main_rtio_core_outputs_record0_seqn2 < main_rtio_core_outputs_record1_seqn2))) begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
		end else begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
		end
		main_rtio_core_outputs_record0_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference0;
		main_rtio_core_outputs_record1_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record0_valid0), main_rtio_core_outputs_record0_payload_channel2} < {(~main_rtio_core_outputs_record1_valid0), main_rtio_core_outputs_record1_payload_channel2})) begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
		end else begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record2_valid0), main_rtio_core_outputs_record2_payload_channel2} == {(~main_rtio_core_outputs_record3_valid0), main_rtio_core_outputs_record3_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record2_seqn2[10] == main_rtio_core_outputs_record2_seqn2[11]) & (main_rtio_core_outputs_record3_seqn2[10] == main_rtio_core_outputs_record3_seqn2[11])) & (main_rtio_core_outputs_record2_seqn2[11] != main_rtio_core_outputs_record3_seqn2[11])) ? main_rtio_core_outputs_record2_seqn2[11] : (main_rtio_core_outputs_record2_seqn2 < main_rtio_core_outputs_record3_seqn2))) begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
		end else begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
		end
		main_rtio_core_outputs_record2_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference1;
		main_rtio_core_outputs_record3_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record2_valid0), main_rtio_core_outputs_record2_payload_channel2} < {(~main_rtio_core_outputs_record3_valid0), main_rtio_core_outputs_record3_payload_channel2})) begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
		end else begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record4_valid0), main_rtio_core_outputs_record4_payload_channel2} == {(~main_rtio_core_outputs_record5_valid0), main_rtio_core_outputs_record5_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record4_seqn2[10] == main_rtio_core_outputs_record4_seqn2[11]) & (main_rtio_core_outputs_record5_seqn2[10] == main_rtio_core_outputs_record5_seqn2[11])) & (main_rtio_core_outputs_record4_seqn2[11] != main_rtio_core_outputs_record5_seqn2[11])) ? main_rtio_core_outputs_record4_seqn2[11] : (main_rtio_core_outputs_record4_seqn2 < main_rtio_core_outputs_record5_seqn2))) begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
		end else begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
		end
		main_rtio_core_outputs_record4_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference2;
		main_rtio_core_outputs_record5_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record4_valid0), main_rtio_core_outputs_record4_payload_channel2} < {(~main_rtio_core_outputs_record5_valid0), main_rtio_core_outputs_record5_payload_channel2})) begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
		end else begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record6_valid0), main_rtio_core_outputs_record6_payload_channel2} == {(~main_rtio_core_outputs_record7_valid0), main_rtio_core_outputs_record7_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record6_seqn2[10] == main_rtio_core_outputs_record6_seqn2[11]) & (main_rtio_core_outputs_record7_seqn2[10] == main_rtio_core_outputs_record7_seqn2[11])) & (main_rtio_core_outputs_record6_seqn2[11] != main_rtio_core_outputs_record7_seqn2[11])) ? main_rtio_core_outputs_record6_seqn2[11] : (main_rtio_core_outputs_record6_seqn2 < main_rtio_core_outputs_record7_seqn2))) begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
		end else begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
		end
		main_rtio_core_outputs_record6_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference3;
		main_rtio_core_outputs_record7_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record6_valid0), main_rtio_core_outputs_record6_payload_channel2} < {(~main_rtio_core_outputs_record7_valid0), main_rtio_core_outputs_record7_payload_channel2})) begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
		end else begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record0_rec_valid), main_rtio_core_outputs_record0_rec_payload_channel} == {(~main_rtio_core_outputs_record2_rec_valid), main_rtio_core_outputs_record2_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record0_rec_seqn[10] == main_rtio_core_outputs_record0_rec_seqn[11]) & (main_rtio_core_outputs_record2_rec_seqn[10] == main_rtio_core_outputs_record2_rec_seqn[11])) & (main_rtio_core_outputs_record0_rec_seqn[11] != main_rtio_core_outputs_record2_rec_seqn[11])) ? main_rtio_core_outputs_record0_rec_seqn[11] : (main_rtio_core_outputs_record0_rec_seqn < main_rtio_core_outputs_record2_rec_seqn))) begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
		end
		main_rtio_core_outputs_record8_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference4;
		main_rtio_core_outputs_record10_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record0_rec_valid), main_rtio_core_outputs_record0_rec_payload_channel} < {(~main_rtio_core_outputs_record2_rec_valid), main_rtio_core_outputs_record2_rec_payload_channel})) begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record1_rec_valid), main_rtio_core_outputs_record1_rec_payload_channel} == {(~main_rtio_core_outputs_record3_rec_valid), main_rtio_core_outputs_record3_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record1_rec_seqn[10] == main_rtio_core_outputs_record1_rec_seqn[11]) & (main_rtio_core_outputs_record3_rec_seqn[10] == main_rtio_core_outputs_record3_rec_seqn[11])) & (main_rtio_core_outputs_record1_rec_seqn[11] != main_rtio_core_outputs_record3_rec_seqn[11])) ? main_rtio_core_outputs_record1_rec_seqn[11] : (main_rtio_core_outputs_record1_rec_seqn < main_rtio_core_outputs_record3_rec_seqn))) begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
		end
		main_rtio_core_outputs_record9_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference5;
		main_rtio_core_outputs_record11_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record1_rec_valid), main_rtio_core_outputs_record1_rec_payload_channel} < {(~main_rtio_core_outputs_record3_rec_valid), main_rtio_core_outputs_record3_rec_payload_channel})) begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record4_rec_valid), main_rtio_core_outputs_record4_rec_payload_channel} == {(~main_rtio_core_outputs_record6_rec_valid), main_rtio_core_outputs_record6_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record4_rec_seqn[10] == main_rtio_core_outputs_record4_rec_seqn[11]) & (main_rtio_core_outputs_record6_rec_seqn[10] == main_rtio_core_outputs_record6_rec_seqn[11])) & (main_rtio_core_outputs_record4_rec_seqn[11] != main_rtio_core_outputs_record6_rec_seqn[11])) ? main_rtio_core_outputs_record4_rec_seqn[11] : (main_rtio_core_outputs_record4_rec_seqn < main_rtio_core_outputs_record6_rec_seqn))) begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
		end
		main_rtio_core_outputs_record12_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference6;
		main_rtio_core_outputs_record14_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record4_rec_valid), main_rtio_core_outputs_record4_rec_payload_channel} < {(~main_rtio_core_outputs_record6_rec_valid), main_rtio_core_outputs_record6_rec_payload_channel})) begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record5_rec_valid), main_rtio_core_outputs_record5_rec_payload_channel} == {(~main_rtio_core_outputs_record7_rec_valid), main_rtio_core_outputs_record7_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record5_rec_seqn[10] == main_rtio_core_outputs_record5_rec_seqn[11]) & (main_rtio_core_outputs_record7_rec_seqn[10] == main_rtio_core_outputs_record7_rec_seqn[11])) & (main_rtio_core_outputs_record5_rec_seqn[11] != main_rtio_core_outputs_record7_rec_seqn[11])) ? main_rtio_core_outputs_record5_rec_seqn[11] : (main_rtio_core_outputs_record5_rec_seqn < main_rtio_core_outputs_record7_rec_seqn))) begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
		end
		main_rtio_core_outputs_record13_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference7;
		main_rtio_core_outputs_record15_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record5_rec_valid), main_rtio_core_outputs_record5_rec_payload_channel} < {(~main_rtio_core_outputs_record7_rec_valid), main_rtio_core_outputs_record7_rec_payload_channel})) begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record9_rec_valid), main_rtio_core_outputs_record9_rec_payload_channel} == {(~main_rtio_core_outputs_record10_rec_valid), main_rtio_core_outputs_record10_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record9_rec_seqn[10] == main_rtio_core_outputs_record9_rec_seqn[11]) & (main_rtio_core_outputs_record10_rec_seqn[10] == main_rtio_core_outputs_record10_rec_seqn[11])) & (main_rtio_core_outputs_record9_rec_seqn[11] != main_rtio_core_outputs_record10_rec_seqn[11])) ? main_rtio_core_outputs_record9_rec_seqn[11] : (main_rtio_core_outputs_record9_rec_seqn < main_rtio_core_outputs_record10_rec_seqn))) begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
		end
		main_rtio_core_outputs_record17_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference8;
		main_rtio_core_outputs_record18_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record9_rec_valid), main_rtio_core_outputs_record9_rec_payload_channel} < {(~main_rtio_core_outputs_record10_rec_valid), main_rtio_core_outputs_record10_rec_payload_channel})) begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record13_rec_valid), main_rtio_core_outputs_record13_rec_payload_channel} == {(~main_rtio_core_outputs_record14_rec_valid), main_rtio_core_outputs_record14_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record13_rec_seqn[10] == main_rtio_core_outputs_record13_rec_seqn[11]) & (main_rtio_core_outputs_record14_rec_seqn[10] == main_rtio_core_outputs_record14_rec_seqn[11])) & (main_rtio_core_outputs_record13_rec_seqn[11] != main_rtio_core_outputs_record14_rec_seqn[11])) ? main_rtio_core_outputs_record13_rec_seqn[11] : (main_rtio_core_outputs_record13_rec_seqn < main_rtio_core_outputs_record14_rec_seqn))) begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
		end
		main_rtio_core_outputs_record21_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference9;
		main_rtio_core_outputs_record22_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record13_rec_valid), main_rtio_core_outputs_record13_rec_payload_channel} < {(~main_rtio_core_outputs_record14_rec_valid), main_rtio_core_outputs_record14_rec_payload_channel})) begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record16_rec_valid <= main_rtio_core_outputs_record8_rec_valid;
	main_rtio_core_outputs_record16_rec_seqn <= main_rtio_core_outputs_record8_rec_seqn;
	main_rtio_core_outputs_record16_rec_replace_occured <= main_rtio_core_outputs_record8_rec_replace_occured;
	main_rtio_core_outputs_record16_rec_nondata_replace_occured <= main_rtio_core_outputs_record8_rec_nondata_replace_occured;
	main_rtio_core_outputs_record16_rec_payload_channel <= main_rtio_core_outputs_record8_rec_payload_channel;
	main_rtio_core_outputs_record16_rec_payload_fine_ts <= main_rtio_core_outputs_record8_rec_payload_fine_ts;
	main_rtio_core_outputs_record16_rec_payload_address <= main_rtio_core_outputs_record8_rec_payload_address;
	main_rtio_core_outputs_record16_rec_payload_data <= main_rtio_core_outputs_record8_rec_payload_data;
	main_rtio_core_outputs_record19_rec_valid <= main_rtio_core_outputs_record11_rec_valid;
	main_rtio_core_outputs_record19_rec_seqn <= main_rtio_core_outputs_record11_rec_seqn;
	main_rtio_core_outputs_record19_rec_replace_occured <= main_rtio_core_outputs_record11_rec_replace_occured;
	main_rtio_core_outputs_record19_rec_nondata_replace_occured <= main_rtio_core_outputs_record11_rec_nondata_replace_occured;
	main_rtio_core_outputs_record19_rec_payload_channel <= main_rtio_core_outputs_record11_rec_payload_channel;
	main_rtio_core_outputs_record19_rec_payload_fine_ts <= main_rtio_core_outputs_record11_rec_payload_fine_ts;
	main_rtio_core_outputs_record19_rec_payload_address <= main_rtio_core_outputs_record11_rec_payload_address;
	main_rtio_core_outputs_record19_rec_payload_data <= main_rtio_core_outputs_record11_rec_payload_data;
	main_rtio_core_outputs_record20_rec_valid <= main_rtio_core_outputs_record12_rec_valid;
	main_rtio_core_outputs_record20_rec_seqn <= main_rtio_core_outputs_record12_rec_seqn;
	main_rtio_core_outputs_record20_rec_replace_occured <= main_rtio_core_outputs_record12_rec_replace_occured;
	main_rtio_core_outputs_record20_rec_nondata_replace_occured <= main_rtio_core_outputs_record12_rec_nondata_replace_occured;
	main_rtio_core_outputs_record20_rec_payload_channel <= main_rtio_core_outputs_record12_rec_payload_channel;
	main_rtio_core_outputs_record20_rec_payload_fine_ts <= main_rtio_core_outputs_record12_rec_payload_fine_ts;
	main_rtio_core_outputs_record20_rec_payload_address <= main_rtio_core_outputs_record12_rec_payload_address;
	main_rtio_core_outputs_record20_rec_payload_data <= main_rtio_core_outputs_record12_rec_payload_data;
	main_rtio_core_outputs_record23_rec_valid <= main_rtio_core_outputs_record15_rec_valid;
	main_rtio_core_outputs_record23_rec_seqn <= main_rtio_core_outputs_record15_rec_seqn;
	main_rtio_core_outputs_record23_rec_replace_occured <= main_rtio_core_outputs_record15_rec_replace_occured;
	main_rtio_core_outputs_record23_rec_nondata_replace_occured <= main_rtio_core_outputs_record15_rec_nondata_replace_occured;
	main_rtio_core_outputs_record23_rec_payload_channel <= main_rtio_core_outputs_record15_rec_payload_channel;
	main_rtio_core_outputs_record23_rec_payload_fine_ts <= main_rtio_core_outputs_record15_rec_payload_fine_ts;
	main_rtio_core_outputs_record23_rec_payload_address <= main_rtio_core_outputs_record15_rec_payload_address;
	main_rtio_core_outputs_record23_rec_payload_data <= main_rtio_core_outputs_record15_rec_payload_data;
	if (({(~main_rtio_core_outputs_record16_rec_valid), main_rtio_core_outputs_record16_rec_payload_channel} == {(~main_rtio_core_outputs_record20_rec_valid), main_rtio_core_outputs_record20_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record16_rec_seqn[10] == main_rtio_core_outputs_record16_rec_seqn[11]) & (main_rtio_core_outputs_record20_rec_seqn[10] == main_rtio_core_outputs_record20_rec_seqn[11])) & (main_rtio_core_outputs_record16_rec_seqn[11] != main_rtio_core_outputs_record20_rec_seqn[11])) ? main_rtio_core_outputs_record16_rec_seqn[11] : (main_rtio_core_outputs_record16_rec_seqn < main_rtio_core_outputs_record20_rec_seqn))) begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
		end
		main_rtio_core_outputs_record24_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference10;
		main_rtio_core_outputs_record28_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record16_rec_valid), main_rtio_core_outputs_record16_rec_payload_channel} < {(~main_rtio_core_outputs_record20_rec_valid), main_rtio_core_outputs_record20_rec_payload_channel})) begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record17_rec_valid), main_rtio_core_outputs_record17_rec_payload_channel} == {(~main_rtio_core_outputs_record21_rec_valid), main_rtio_core_outputs_record21_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record17_rec_seqn[10] == main_rtio_core_outputs_record17_rec_seqn[11]) & (main_rtio_core_outputs_record21_rec_seqn[10] == main_rtio_core_outputs_record21_rec_seqn[11])) & (main_rtio_core_outputs_record17_rec_seqn[11] != main_rtio_core_outputs_record21_rec_seqn[11])) ? main_rtio_core_outputs_record17_rec_seqn[11] : (main_rtio_core_outputs_record17_rec_seqn < main_rtio_core_outputs_record21_rec_seqn))) begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
		end
		main_rtio_core_outputs_record25_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference11;
		main_rtio_core_outputs_record29_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record17_rec_valid), main_rtio_core_outputs_record17_rec_payload_channel} < {(~main_rtio_core_outputs_record21_rec_valid), main_rtio_core_outputs_record21_rec_payload_channel})) begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record18_rec_valid), main_rtio_core_outputs_record18_rec_payload_channel} == {(~main_rtio_core_outputs_record22_rec_valid), main_rtio_core_outputs_record22_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record18_rec_seqn[10] == main_rtio_core_outputs_record18_rec_seqn[11]) & (main_rtio_core_outputs_record22_rec_seqn[10] == main_rtio_core_outputs_record22_rec_seqn[11])) & (main_rtio_core_outputs_record18_rec_seqn[11] != main_rtio_core_outputs_record22_rec_seqn[11])) ? main_rtio_core_outputs_record18_rec_seqn[11] : (main_rtio_core_outputs_record18_rec_seqn < main_rtio_core_outputs_record22_rec_seqn))) begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
		end
		main_rtio_core_outputs_record26_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference12;
		main_rtio_core_outputs_record30_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record18_rec_valid), main_rtio_core_outputs_record18_rec_payload_channel} < {(~main_rtio_core_outputs_record22_rec_valid), main_rtio_core_outputs_record22_rec_payload_channel})) begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record19_rec_valid), main_rtio_core_outputs_record19_rec_payload_channel} == {(~main_rtio_core_outputs_record23_rec_valid), main_rtio_core_outputs_record23_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record19_rec_seqn[10] == main_rtio_core_outputs_record19_rec_seqn[11]) & (main_rtio_core_outputs_record23_rec_seqn[10] == main_rtio_core_outputs_record23_rec_seqn[11])) & (main_rtio_core_outputs_record19_rec_seqn[11] != main_rtio_core_outputs_record23_rec_seqn[11])) ? main_rtio_core_outputs_record19_rec_seqn[11] : (main_rtio_core_outputs_record19_rec_seqn < main_rtio_core_outputs_record23_rec_seqn))) begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
		end
		main_rtio_core_outputs_record27_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference13;
		main_rtio_core_outputs_record31_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record19_rec_valid), main_rtio_core_outputs_record19_rec_payload_channel} < {(~main_rtio_core_outputs_record23_rec_valid), main_rtio_core_outputs_record23_rec_payload_channel})) begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record26_rec_valid), main_rtio_core_outputs_record26_rec_payload_channel} == {(~main_rtio_core_outputs_record28_rec_valid), main_rtio_core_outputs_record28_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record26_rec_seqn[10] == main_rtio_core_outputs_record26_rec_seqn[11]) & (main_rtio_core_outputs_record28_rec_seqn[10] == main_rtio_core_outputs_record28_rec_seqn[11])) & (main_rtio_core_outputs_record26_rec_seqn[11] != main_rtio_core_outputs_record28_rec_seqn[11])) ? main_rtio_core_outputs_record26_rec_seqn[11] : (main_rtio_core_outputs_record26_rec_seqn < main_rtio_core_outputs_record28_rec_seqn))) begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
		end
		main_rtio_core_outputs_record34_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference14;
		main_rtio_core_outputs_record36_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record26_rec_valid), main_rtio_core_outputs_record26_rec_payload_channel} < {(~main_rtio_core_outputs_record28_rec_valid), main_rtio_core_outputs_record28_rec_payload_channel})) begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record27_rec_valid), main_rtio_core_outputs_record27_rec_payload_channel} == {(~main_rtio_core_outputs_record29_rec_valid), main_rtio_core_outputs_record29_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record27_rec_seqn[10] == main_rtio_core_outputs_record27_rec_seqn[11]) & (main_rtio_core_outputs_record29_rec_seqn[10] == main_rtio_core_outputs_record29_rec_seqn[11])) & (main_rtio_core_outputs_record27_rec_seqn[11] != main_rtio_core_outputs_record29_rec_seqn[11])) ? main_rtio_core_outputs_record27_rec_seqn[11] : (main_rtio_core_outputs_record27_rec_seqn < main_rtio_core_outputs_record29_rec_seqn))) begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
		end
		main_rtio_core_outputs_record35_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference15;
		main_rtio_core_outputs_record37_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record27_rec_valid), main_rtio_core_outputs_record27_rec_payload_channel} < {(~main_rtio_core_outputs_record29_rec_valid), main_rtio_core_outputs_record29_rec_payload_channel})) begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record32_rec_valid <= main_rtio_core_outputs_record24_rec_valid;
	main_rtio_core_outputs_record32_rec_seqn <= main_rtio_core_outputs_record24_rec_seqn;
	main_rtio_core_outputs_record32_rec_replace_occured <= main_rtio_core_outputs_record24_rec_replace_occured;
	main_rtio_core_outputs_record32_rec_nondata_replace_occured <= main_rtio_core_outputs_record24_rec_nondata_replace_occured;
	main_rtio_core_outputs_record32_rec_payload_channel <= main_rtio_core_outputs_record24_rec_payload_channel;
	main_rtio_core_outputs_record32_rec_payload_fine_ts <= main_rtio_core_outputs_record24_rec_payload_fine_ts;
	main_rtio_core_outputs_record32_rec_payload_address <= main_rtio_core_outputs_record24_rec_payload_address;
	main_rtio_core_outputs_record32_rec_payload_data <= main_rtio_core_outputs_record24_rec_payload_data;
	main_rtio_core_outputs_record33_rec_valid <= main_rtio_core_outputs_record25_rec_valid;
	main_rtio_core_outputs_record33_rec_seqn <= main_rtio_core_outputs_record25_rec_seqn;
	main_rtio_core_outputs_record33_rec_replace_occured <= main_rtio_core_outputs_record25_rec_replace_occured;
	main_rtio_core_outputs_record33_rec_nondata_replace_occured <= main_rtio_core_outputs_record25_rec_nondata_replace_occured;
	main_rtio_core_outputs_record33_rec_payload_channel <= main_rtio_core_outputs_record25_rec_payload_channel;
	main_rtio_core_outputs_record33_rec_payload_fine_ts <= main_rtio_core_outputs_record25_rec_payload_fine_ts;
	main_rtio_core_outputs_record33_rec_payload_address <= main_rtio_core_outputs_record25_rec_payload_address;
	main_rtio_core_outputs_record33_rec_payload_data <= main_rtio_core_outputs_record25_rec_payload_data;
	main_rtio_core_outputs_record38_rec_valid <= main_rtio_core_outputs_record30_rec_valid;
	main_rtio_core_outputs_record38_rec_seqn <= main_rtio_core_outputs_record30_rec_seqn;
	main_rtio_core_outputs_record38_rec_replace_occured <= main_rtio_core_outputs_record30_rec_replace_occured;
	main_rtio_core_outputs_record38_rec_nondata_replace_occured <= main_rtio_core_outputs_record30_rec_nondata_replace_occured;
	main_rtio_core_outputs_record38_rec_payload_channel <= main_rtio_core_outputs_record30_rec_payload_channel;
	main_rtio_core_outputs_record38_rec_payload_fine_ts <= main_rtio_core_outputs_record30_rec_payload_fine_ts;
	main_rtio_core_outputs_record38_rec_payload_address <= main_rtio_core_outputs_record30_rec_payload_address;
	main_rtio_core_outputs_record38_rec_payload_data <= main_rtio_core_outputs_record30_rec_payload_data;
	main_rtio_core_outputs_record39_rec_valid <= main_rtio_core_outputs_record31_rec_valid;
	main_rtio_core_outputs_record39_rec_seqn <= main_rtio_core_outputs_record31_rec_seqn;
	main_rtio_core_outputs_record39_rec_replace_occured <= main_rtio_core_outputs_record31_rec_replace_occured;
	main_rtio_core_outputs_record39_rec_nondata_replace_occured <= main_rtio_core_outputs_record31_rec_nondata_replace_occured;
	main_rtio_core_outputs_record39_rec_payload_channel <= main_rtio_core_outputs_record31_rec_payload_channel;
	main_rtio_core_outputs_record39_rec_payload_fine_ts <= main_rtio_core_outputs_record31_rec_payload_fine_ts;
	main_rtio_core_outputs_record39_rec_payload_address <= main_rtio_core_outputs_record31_rec_payload_address;
	main_rtio_core_outputs_record39_rec_payload_data <= main_rtio_core_outputs_record31_rec_payload_data;
	if (({(~main_rtio_core_outputs_record33_rec_valid), main_rtio_core_outputs_record33_rec_payload_channel} == {(~main_rtio_core_outputs_record34_rec_valid), main_rtio_core_outputs_record34_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record33_rec_seqn[10] == main_rtio_core_outputs_record33_rec_seqn[11]) & (main_rtio_core_outputs_record34_rec_seqn[10] == main_rtio_core_outputs_record34_rec_seqn[11])) & (main_rtio_core_outputs_record33_rec_seqn[11] != main_rtio_core_outputs_record34_rec_seqn[11])) ? main_rtio_core_outputs_record33_rec_seqn[11] : (main_rtio_core_outputs_record33_rec_seqn < main_rtio_core_outputs_record34_rec_seqn))) begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
		end
		main_rtio_core_outputs_record41_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference16;
		main_rtio_core_outputs_record42_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record33_rec_valid), main_rtio_core_outputs_record33_rec_payload_channel} < {(~main_rtio_core_outputs_record34_rec_valid), main_rtio_core_outputs_record34_rec_payload_channel})) begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record35_rec_valid), main_rtio_core_outputs_record35_rec_payload_channel} == {(~main_rtio_core_outputs_record36_rec_valid), main_rtio_core_outputs_record36_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record35_rec_seqn[10] == main_rtio_core_outputs_record35_rec_seqn[11]) & (main_rtio_core_outputs_record36_rec_seqn[10] == main_rtio_core_outputs_record36_rec_seqn[11])) & (main_rtio_core_outputs_record35_rec_seqn[11] != main_rtio_core_outputs_record36_rec_seqn[11])) ? main_rtio_core_outputs_record35_rec_seqn[11] : (main_rtio_core_outputs_record35_rec_seqn < main_rtio_core_outputs_record36_rec_seqn))) begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
		end
		main_rtio_core_outputs_record43_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference17;
		main_rtio_core_outputs_record44_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record35_rec_valid), main_rtio_core_outputs_record35_rec_payload_channel} < {(~main_rtio_core_outputs_record36_rec_valid), main_rtio_core_outputs_record36_rec_payload_channel})) begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record37_rec_valid), main_rtio_core_outputs_record37_rec_payload_channel} == {(~main_rtio_core_outputs_record38_rec_valid), main_rtio_core_outputs_record38_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record37_rec_seqn[10] == main_rtio_core_outputs_record37_rec_seqn[11]) & (main_rtio_core_outputs_record38_rec_seqn[10] == main_rtio_core_outputs_record38_rec_seqn[11])) & (main_rtio_core_outputs_record37_rec_seqn[11] != main_rtio_core_outputs_record38_rec_seqn[11])) ? main_rtio_core_outputs_record37_rec_seqn[11] : (main_rtio_core_outputs_record37_rec_seqn < main_rtio_core_outputs_record38_rec_seqn))) begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
		end
		main_rtio_core_outputs_record45_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference18;
		main_rtio_core_outputs_record46_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record37_rec_valid), main_rtio_core_outputs_record37_rec_payload_channel} < {(~main_rtio_core_outputs_record38_rec_valid), main_rtio_core_outputs_record38_rec_payload_channel})) begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record40_rec_valid <= main_rtio_core_outputs_record32_rec_valid;
	main_rtio_core_outputs_record40_rec_seqn <= main_rtio_core_outputs_record32_rec_seqn;
	main_rtio_core_outputs_record40_rec_replace_occured <= main_rtio_core_outputs_record32_rec_replace_occured;
	main_rtio_core_outputs_record40_rec_nondata_replace_occured <= main_rtio_core_outputs_record32_rec_nondata_replace_occured;
	main_rtio_core_outputs_record40_rec_payload_channel <= main_rtio_core_outputs_record32_rec_payload_channel;
	main_rtio_core_outputs_record40_rec_payload_fine_ts <= main_rtio_core_outputs_record32_rec_payload_fine_ts;
	main_rtio_core_outputs_record40_rec_payload_address <= main_rtio_core_outputs_record32_rec_payload_address;
	main_rtio_core_outputs_record40_rec_payload_data <= main_rtio_core_outputs_record32_rec_payload_data;
	main_rtio_core_outputs_record47_rec_valid <= main_rtio_core_outputs_record39_rec_valid;
	main_rtio_core_outputs_record47_rec_seqn <= main_rtio_core_outputs_record39_rec_seqn;
	main_rtio_core_outputs_record47_rec_replace_occured <= main_rtio_core_outputs_record39_rec_replace_occured;
	main_rtio_core_outputs_record47_rec_nondata_replace_occured <= main_rtio_core_outputs_record39_rec_nondata_replace_occured;
	main_rtio_core_outputs_record47_rec_payload_channel <= main_rtio_core_outputs_record39_rec_payload_channel;
	main_rtio_core_outputs_record47_rec_payload_fine_ts <= main_rtio_core_outputs_record39_rec_payload_fine_ts;
	main_rtio_core_outputs_record47_rec_payload_address <= main_rtio_core_outputs_record39_rec_payload_address;
	main_rtio_core_outputs_record47_rec_payload_data <= main_rtio_core_outputs_record39_rec_payload_data;
	main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
	main_rtio_core_inputs_asyncfifo0_graycounter0_q <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
	if (main_rtio_core_inputs_blindtransfer0_i) begin
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer0_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer0_ps_i) begin
		main_rtio_core_inputs_blindtransfer0_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer0_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
	main_rtio_core_inputs_asyncfifo1_graycounter2_q <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
	if (main_rtio_core_inputs_blindtransfer1_i) begin
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer1_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer1_ps_i) begin
		main_rtio_core_inputs_blindtransfer1_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer1_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
	main_rtio_core_inputs_asyncfifo2_graycounter4_q <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
	if (main_rtio_core_inputs_blindtransfer2_i) begin
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer2_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer2_ps_i) begin
		main_rtio_core_inputs_blindtransfer2_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer2_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
	main_rtio_core_inputs_asyncfifo3_graycounter6_q <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
	if (main_rtio_core_inputs_blindtransfer3_i) begin
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer3_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer3_ps_i) begin
		main_rtio_core_inputs_blindtransfer3_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer3_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
	main_rtio_core_inputs_asyncfifo4_graycounter8_q <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
	if (main_rtio_core_inputs_blindtransfer4_i) begin
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer4_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer4_ps_i) begin
		main_rtio_core_inputs_blindtransfer4_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer4_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
	main_rtio_core_inputs_asyncfifo5_graycounter10_q <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
	if (main_rtio_core_inputs_blindtransfer5_i) begin
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer5_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer5_ps_i) begin
		main_rtio_core_inputs_blindtransfer5_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer5_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
	main_rtio_core_inputs_asyncfifo6_graycounter12_q <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
	if (main_rtio_core_inputs_blindtransfer6_i) begin
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer6_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer6_ps_i) begin
		main_rtio_core_inputs_blindtransfer6_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer6_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary;
	main_rtio_core_inputs_asyncfifo7_graycounter14_q <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_next;
	if (main_rtio_core_inputs_blindtransfer7_i) begin
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer7_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer7_ps_i) begin
		main_rtio_core_inputs_blindtransfer7_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer7_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary;
	main_rtio_core_inputs_asyncfifo8_graycounter16_q <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_next;
	if (main_rtio_core_inputs_blindtransfer8_i) begin
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer8_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer8_ps_i) begin
		main_rtio_core_inputs_blindtransfer8_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer8_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary;
	main_rtio_core_inputs_asyncfifo9_graycounter18_q <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_next;
	if (main_rtio_core_inputs_blindtransfer9_i) begin
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer9_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer9_ps_i) begin
		main_rtio_core_inputs_blindtransfer9_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer9_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary;
	main_rtio_core_inputs_asyncfifo10_graycounter20_q <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_next;
	if (main_rtio_core_inputs_blindtransfer10_i) begin
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer10_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer10_ps_i) begin
		main_rtio_core_inputs_blindtransfer10_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer10_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o;
	if (main_rtio_core_o_collision_sync_i) begin
		main_rtio_core_o_collision_sync_blind <= 1'd1;
	end
	if (main_rtio_core_o_collision_sync_ps_ack_o) begin
		main_rtio_core_o_collision_sync_blind <= 1'd0;
	end
	if (main_rtio_core_o_collision_sync_ps_i) begin
		main_rtio_core_o_collision_sync_bxfer_data <= main_rtio_core_o_collision_sync_data_i;
	end
	if (main_rtio_core_o_collision_sync_ps_i) begin
		main_rtio_core_o_collision_sync_ps_toggle_i <= (~main_rtio_core_o_collision_sync_ps_toggle_i);
	end
	main_rtio_core_o_collision_sync_ps_ack_toggle_o_r <= main_rtio_core_o_collision_sync_ps_ack_toggle_o;
	if (main_rtio_core_o_busy_sync_i) begin
		main_rtio_core_o_busy_sync_blind <= 1'd1;
	end
	if (main_rtio_core_o_busy_sync_ps_ack_o) begin
		main_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	if (main_rtio_core_o_busy_sync_ps_i) begin
		main_rtio_core_o_busy_sync_bxfer_data <= main_rtio_core_o_busy_sync_data_i;
	end
	if (main_rtio_core_o_busy_sync_ps_i) begin
		main_rtio_core_o_busy_sync_ps_toggle_i <= (~main_rtio_core_o_busy_sync_ps_toggle_i);
	end
	main_rtio_core_o_busy_sync_ps_ack_toggle_o_r <= main_rtio_core_o_busy_sync_ps_ack_toggle_o;
	if (rio_rst) begin
		main_inout_8x0_inout_8x0_ointerface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_sensitivity <= 2'd0;
		main_inout_8x0_inout_8x0_sample <= 1'd0;
		main_inout_8x1_inout_8x1_ointerface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_sensitivity <= 2'd0;
		main_inout_8x1_inout_8x1_sample <= 1'd0;
		main_inout_8x2_inout_8x2_ointerface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_sensitivity <= 2'd0;
		main_inout_8x2_inout_8x2_sample <= 1'd0;
		main_inout_8x3_inout_8x3_ointerface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_sensitivity <= 2'd0;
		main_inout_8x3_inout_8x3_sample <= 1'd0;
		main_inout_8x4_inout_8x4_ointerface4_stb <= 1'd0;
		main_inout_8x4_inout_8x4_sensitivity <= 2'd0;
		main_inout_8x4_inout_8x4_sample <= 1'd0;
		main_inout_8x5_inout_8x5_ointerface5_stb <= 1'd0;
		main_inout_8x5_inout_8x5_sensitivity <= 2'd0;
		main_inout_8x5_inout_8x5_sample <= 1'd0;
		main_inout_8x6_inout_8x6_ointerface6_stb <= 1'd0;
		main_inout_8x6_inout_8x6_sensitivity <= 2'd0;
		main_inout_8x6_inout_8x6_sample <= 1'd0;
		main_inout_8x7_inout_8x7_ointerface7_stb <= 1'd0;
		main_inout_8x7_inout_8x7_sensitivity <= 2'd0;
		main_inout_8x7_inout_8x7_sample <= 1'd0;
		main_output_8x0_stb <= 1'd0;
		main_output_8x1_stb <= 1'd0;
		main_output_8x2_stb <= 1'd0;
		main_output_8x3_stb <= 1'd0;
		main_output_8x4_stb <= 1'd0;
		main_output_8x5_stb <= 1'd0;
		main_output_8x6_stb <= 1'd0;
		main_output_8x7_stb <= 1'd0;
		main_spimaster0_ointerface0_stb <= 1'd0;
		main_output_8x8_stb <= 1'd0;
		main_output_8x9_stb <= 1'd0;
		main_output_8x10_stb <= 1'd0;
		main_output_8x11_stb <= 1'd0;
		main_output_8x12_stb <= 1'd0;
		main_spimaster1_ointerface1_stb <= 1'd0;
		main_output_8x13_stb <= 1'd0;
		main_output_8x14_stb <= 1'd0;
		main_output_8x15_stb <= 1'd0;
		main_output_8x16_stb <= 1'd0;
		main_output_8x17_stb <= 1'd0;
		main_spimaster2_ointerface2_stb <= 1'd0;
		main_output_8x18_stb <= 1'd0;
		main_output_8x19_stb <= 1'd0;
		main_output_8x20_stb <= 1'd0;
		main_output_8x21_stb <= 1'd0;
		main_output_8x22_stb <= 1'd0;
		main_output0_stb <= 1'd0;
		main_output1_stb <= 1'd0;
		main_stb <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered0_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= 8'd0;
		main_rtio_core_outputs_gates_record0_valid <= 1'd0;
		main_rtio_core_outputs_gates_record1_valid <= 1'd0;
		main_rtio_core_outputs_gates_record2_valid <= 1'd0;
		main_rtio_core_outputs_gates_record3_valid <= 1'd0;
		main_rtio_core_outputs_gates_record4_valid <= 1'd0;
		main_rtio_core_outputs_gates_record5_valid <= 1'd0;
		main_rtio_core_outputs_gates_record6_valid <= 1'd0;
		main_rtio_core_outputs_gates_record7_valid <= 1'd0;
		main_rtio_core_outputs_collision <= 1'd0;
		main_rtio_core_outputs_busy <= 1'd0;
		main_rtio_core_outputs_record0_rec_valid <= 1'd0;
		main_rtio_core_outputs_record1_rec_valid <= 1'd0;
		main_rtio_core_outputs_record2_rec_valid <= 1'd0;
		main_rtio_core_outputs_record3_rec_valid <= 1'd0;
		main_rtio_core_outputs_record4_rec_valid <= 1'd0;
		main_rtio_core_outputs_record5_rec_valid <= 1'd0;
		main_rtio_core_outputs_record6_rec_valid <= 1'd0;
		main_rtio_core_outputs_record7_rec_valid <= 1'd0;
		main_rtio_core_outputs_record8_rec_valid <= 1'd0;
		main_rtio_core_outputs_record9_rec_valid <= 1'd0;
		main_rtio_core_outputs_record10_rec_valid <= 1'd0;
		main_rtio_core_outputs_record11_rec_valid <= 1'd0;
		main_rtio_core_outputs_record12_rec_valid <= 1'd0;
		main_rtio_core_outputs_record13_rec_valid <= 1'd0;
		main_rtio_core_outputs_record14_rec_valid <= 1'd0;
		main_rtio_core_outputs_record15_rec_valid <= 1'd0;
		main_rtio_core_outputs_record16_rec_valid <= 1'd0;
		main_rtio_core_outputs_record17_rec_valid <= 1'd0;
		main_rtio_core_outputs_record18_rec_valid <= 1'd0;
		main_rtio_core_outputs_record19_rec_valid <= 1'd0;
		main_rtio_core_outputs_record20_rec_valid <= 1'd0;
		main_rtio_core_outputs_record21_rec_valid <= 1'd0;
		main_rtio_core_outputs_record22_rec_valid <= 1'd0;
		main_rtio_core_outputs_record23_rec_valid <= 1'd0;
		main_rtio_core_outputs_record24_rec_valid <= 1'd0;
		main_rtio_core_outputs_record25_rec_valid <= 1'd0;
		main_rtio_core_outputs_record26_rec_valid <= 1'd0;
		main_rtio_core_outputs_record27_rec_valid <= 1'd0;
		main_rtio_core_outputs_record28_rec_valid <= 1'd0;
		main_rtio_core_outputs_record29_rec_valid <= 1'd0;
		main_rtio_core_outputs_record30_rec_valid <= 1'd0;
		main_rtio_core_outputs_record31_rec_valid <= 1'd0;
		main_rtio_core_outputs_record32_rec_valid <= 1'd0;
		main_rtio_core_outputs_record33_rec_valid <= 1'd0;
		main_rtio_core_outputs_record34_rec_valid <= 1'd0;
		main_rtio_core_outputs_record35_rec_valid <= 1'd0;
		main_rtio_core_outputs_record36_rec_valid <= 1'd0;
		main_rtio_core_outputs_record37_rec_valid <= 1'd0;
		main_rtio_core_outputs_record38_rec_valid <= 1'd0;
		main_rtio_core_outputs_record39_rec_valid <= 1'd0;
		main_rtio_core_outputs_record40_rec_valid <= 1'd0;
		main_rtio_core_outputs_record41_rec_valid <= 1'd0;
		main_rtio_core_outputs_record42_rec_valid <= 1'd0;
		main_rtio_core_outputs_record43_rec_valid <= 1'd0;
		main_rtio_core_outputs_record44_rec_valid <= 1'd0;
		main_rtio_core_outputs_record45_rec_valid <= 1'd0;
		main_rtio_core_outputs_record46_rec_valid <= 1'd0;
		main_rtio_core_outputs_record47_rec_valid <= 1'd0;
		main_rtio_core_outputs_record0_valid1 <= 1'd0;
		main_rtio_core_outputs_record1_valid1 <= 1'd0;
		main_rtio_core_outputs_record2_valid1 <= 1'd0;
		main_rtio_core_outputs_record3_valid1 <= 1'd0;
		main_rtio_core_outputs_record4_valid1 <= 1'd0;
		main_rtio_core_outputs_record5_valid1 <= 1'd0;
		main_rtio_core_outputs_record6_valid1 <= 1'd0;
		main_rtio_core_outputs_record7_valid1 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r0 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r0 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r1 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r1 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r2 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r2 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r3 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r3 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r4 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r4 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r5 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r5 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r6 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r6 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r7 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r7 <= 1'd0;
		main_rtio_core_outputs_stb_r0 <= 1'd0;
		main_rtio_core_outputs_stb_r1 <= 1'd0;
		main_rtio_core_outputs_stb_r2 <= 1'd0;
		main_rtio_core_outputs_stb_r3 <= 1'd0;
		main_rtio_core_outputs_stb_r4 <= 1'd0;
		main_rtio_core_outputs_stb_r5 <= 1'd0;
		main_rtio_core_outputs_stb_r6 <= 1'd0;
		main_rtio_core_outputs_stb_r7 <= 1'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter0_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter2_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter4_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter6_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter8_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter10_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter12_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter14_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary <= 7'd0;
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter16_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary <= 3'd0;
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter18_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary <= 3'd0;
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter20_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary <= 3'd0;
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd0;
		main_rtio_core_o_collision_sync_blind <= 1'd0;
		main_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	builder_xilinxmultiregimpl17_regs0 <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q;
	builder_xilinxmultiregimpl17_regs1 <= builder_xilinxmultiregimpl17_regs0;
	builder_xilinxmultiregimpl19_regs0 <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q;
	builder_xilinxmultiregimpl19_regs1 <= builder_xilinxmultiregimpl19_regs0;
	builder_xilinxmultiregimpl21_regs0 <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q;
	builder_xilinxmultiregimpl21_regs1 <= builder_xilinxmultiregimpl21_regs0;
	builder_xilinxmultiregimpl23_regs0 <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q;
	builder_xilinxmultiregimpl23_regs1 <= builder_xilinxmultiregimpl23_regs0;
	builder_xilinxmultiregimpl25_regs0 <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q;
	builder_xilinxmultiregimpl25_regs1 <= builder_xilinxmultiregimpl25_regs0;
	builder_xilinxmultiregimpl27_regs0 <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q;
	builder_xilinxmultiregimpl27_regs1 <= builder_xilinxmultiregimpl27_regs0;
	builder_xilinxmultiregimpl29_regs0 <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q;
	builder_xilinxmultiregimpl29_regs1 <= builder_xilinxmultiregimpl29_regs0;
	builder_xilinxmultiregimpl31_regs0 <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q;
	builder_xilinxmultiregimpl31_regs1 <= builder_xilinxmultiregimpl31_regs0;
	builder_xilinxmultiregimpl34_regs0 <= main_rtio_core_inputs_asyncfifo0_graycounter1_q;
	builder_xilinxmultiregimpl34_regs1 <= builder_xilinxmultiregimpl34_regs0;
	builder_xilinxmultiregimpl36_regs0 <= main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i;
	builder_xilinxmultiregimpl36_regs1 <= builder_xilinxmultiregimpl36_regs0;
	builder_xilinxmultiregimpl38_regs0 <= main_rtio_core_inputs_asyncfifo1_graycounter3_q;
	builder_xilinxmultiregimpl38_regs1 <= builder_xilinxmultiregimpl38_regs0;
	builder_xilinxmultiregimpl40_regs0 <= main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i;
	builder_xilinxmultiregimpl40_regs1 <= builder_xilinxmultiregimpl40_regs0;
	builder_xilinxmultiregimpl42_regs0 <= main_rtio_core_inputs_asyncfifo2_graycounter5_q;
	builder_xilinxmultiregimpl42_regs1 <= builder_xilinxmultiregimpl42_regs0;
	builder_xilinxmultiregimpl44_regs0 <= main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i;
	builder_xilinxmultiregimpl44_regs1 <= builder_xilinxmultiregimpl44_regs0;
	builder_xilinxmultiregimpl46_regs0 <= main_rtio_core_inputs_asyncfifo3_graycounter7_q;
	builder_xilinxmultiregimpl46_regs1 <= builder_xilinxmultiregimpl46_regs0;
	builder_xilinxmultiregimpl48_regs0 <= main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i;
	builder_xilinxmultiregimpl48_regs1 <= builder_xilinxmultiregimpl48_regs0;
	builder_xilinxmultiregimpl50_regs0 <= main_rtio_core_inputs_asyncfifo4_graycounter9_q;
	builder_xilinxmultiregimpl50_regs1 <= builder_xilinxmultiregimpl50_regs0;
	builder_xilinxmultiregimpl52_regs0 <= main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i;
	builder_xilinxmultiregimpl52_regs1 <= builder_xilinxmultiregimpl52_regs0;
	builder_xilinxmultiregimpl54_regs0 <= main_rtio_core_inputs_asyncfifo5_graycounter11_q;
	builder_xilinxmultiregimpl54_regs1 <= builder_xilinxmultiregimpl54_regs0;
	builder_xilinxmultiregimpl56_regs0 <= main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i;
	builder_xilinxmultiregimpl56_regs1 <= builder_xilinxmultiregimpl56_regs0;
	builder_xilinxmultiregimpl58_regs0 <= main_rtio_core_inputs_asyncfifo6_graycounter13_q;
	builder_xilinxmultiregimpl58_regs1 <= builder_xilinxmultiregimpl58_regs0;
	builder_xilinxmultiregimpl60_regs0 <= main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i;
	builder_xilinxmultiregimpl60_regs1 <= builder_xilinxmultiregimpl60_regs0;
	builder_xilinxmultiregimpl62_regs0 <= main_rtio_core_inputs_asyncfifo7_graycounter15_q;
	builder_xilinxmultiregimpl62_regs1 <= builder_xilinxmultiregimpl62_regs0;
	builder_xilinxmultiregimpl64_regs0 <= main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i;
	builder_xilinxmultiregimpl64_regs1 <= builder_xilinxmultiregimpl64_regs0;
	builder_xilinxmultiregimpl66_regs0 <= main_rtio_core_inputs_asyncfifo8_graycounter17_q;
	builder_xilinxmultiregimpl66_regs1 <= builder_xilinxmultiregimpl66_regs0;
	builder_xilinxmultiregimpl68_regs0 <= main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i;
	builder_xilinxmultiregimpl68_regs1 <= builder_xilinxmultiregimpl68_regs0;
	builder_xilinxmultiregimpl70_regs0 <= main_rtio_core_inputs_asyncfifo9_graycounter19_q;
	builder_xilinxmultiregimpl70_regs1 <= builder_xilinxmultiregimpl70_regs0;
	builder_xilinxmultiregimpl72_regs0 <= main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i;
	builder_xilinxmultiregimpl72_regs1 <= builder_xilinxmultiregimpl72_regs0;
	builder_xilinxmultiregimpl74_regs0 <= main_rtio_core_inputs_asyncfifo10_graycounter21_q;
	builder_xilinxmultiregimpl74_regs1 <= builder_xilinxmultiregimpl74_regs0;
	builder_xilinxmultiregimpl76_regs0 <= main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i;
	builder_xilinxmultiregimpl76_regs1 <= builder_xilinxmultiregimpl76_regs0;
	builder_xilinxmultiregimpl78_regs0 <= main_rtio_core_o_collision_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl78_regs1 <= builder_xilinxmultiregimpl78_regs0;
	builder_xilinxmultiregimpl81_regs0 <= main_rtio_core_o_busy_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl81_regs1 <= builder_xilinxmultiregimpl81_regs0;
	builder_xilinxmultiregimpl124_regs0 <= main_inj_o_sys0;
	builder_xilinxmultiregimpl124_regs1 <= builder_xilinxmultiregimpl124_regs0;
	builder_xilinxmultiregimpl125_regs0 <= main_inj_o_sys1;
	builder_xilinxmultiregimpl125_regs1 <= builder_xilinxmultiregimpl125_regs0;
	builder_xilinxmultiregimpl126_regs0 <= main_inj_o_sys2;
	builder_xilinxmultiregimpl126_regs1 <= builder_xilinxmultiregimpl126_regs0;
	builder_xilinxmultiregimpl127_regs0 <= main_inj_o_sys3;
	builder_xilinxmultiregimpl127_regs1 <= builder_xilinxmultiregimpl127_regs0;
	builder_xilinxmultiregimpl128_regs0 <= main_inj_o_sys4;
	builder_xilinxmultiregimpl128_regs1 <= builder_xilinxmultiregimpl128_regs0;
	builder_xilinxmultiregimpl129_regs0 <= main_inj_o_sys5;
	builder_xilinxmultiregimpl129_regs1 <= builder_xilinxmultiregimpl129_regs0;
	builder_xilinxmultiregimpl130_regs0 <= main_inj_o_sys6;
	builder_xilinxmultiregimpl130_regs1 <= builder_xilinxmultiregimpl130_regs0;
	builder_xilinxmultiregimpl131_regs0 <= main_inj_o_sys7;
	builder_xilinxmultiregimpl131_regs1 <= builder_xilinxmultiregimpl131_regs0;
	builder_xilinxmultiregimpl132_regs0 <= main_inj_o_sys8;
	builder_xilinxmultiregimpl132_regs1 <= builder_xilinxmultiregimpl132_regs0;
	builder_xilinxmultiregimpl133_regs0 <= main_inj_o_sys9;
	builder_xilinxmultiregimpl133_regs1 <= builder_xilinxmultiregimpl133_regs0;
	builder_xilinxmultiregimpl134_regs0 <= main_inj_o_sys10;
	builder_xilinxmultiregimpl134_regs1 <= builder_xilinxmultiregimpl134_regs0;
	builder_xilinxmultiregimpl135_regs0 <= main_inj_o_sys11;
	builder_xilinxmultiregimpl135_regs1 <= builder_xilinxmultiregimpl135_regs0;
	builder_xilinxmultiregimpl136_regs0 <= main_inj_o_sys12;
	builder_xilinxmultiregimpl136_regs1 <= builder_xilinxmultiregimpl136_regs0;
	builder_xilinxmultiregimpl137_regs0 <= main_inj_o_sys13;
	builder_xilinxmultiregimpl137_regs1 <= builder_xilinxmultiregimpl137_regs0;
	builder_xilinxmultiregimpl138_regs0 <= main_inj_o_sys14;
	builder_xilinxmultiregimpl138_regs1 <= builder_xilinxmultiregimpl138_regs0;
	builder_xilinxmultiregimpl139_regs0 <= main_inj_o_sys15;
	builder_xilinxmultiregimpl139_regs1 <= builder_xilinxmultiregimpl139_regs0;
	builder_xilinxmultiregimpl140_regs0 <= main_inj_o_sys16;
	builder_xilinxmultiregimpl140_regs1 <= builder_xilinxmultiregimpl140_regs0;
	builder_xilinxmultiregimpl141_regs0 <= main_inj_o_sys17;
	builder_xilinxmultiregimpl141_regs1 <= builder_xilinxmultiregimpl141_regs0;
	builder_xilinxmultiregimpl142_regs0 <= main_inj_o_sys18;
	builder_xilinxmultiregimpl142_regs1 <= builder_xilinxmultiregimpl142_regs0;
	builder_xilinxmultiregimpl143_regs0 <= main_inj_o_sys19;
	builder_xilinxmultiregimpl143_regs1 <= builder_xilinxmultiregimpl143_regs0;
	builder_xilinxmultiregimpl144_regs0 <= main_inj_o_sys20;
	builder_xilinxmultiregimpl144_regs1 <= builder_xilinxmultiregimpl144_regs0;
	builder_xilinxmultiregimpl145_regs0 <= main_inj_o_sys21;
	builder_xilinxmultiregimpl145_regs1 <= builder_xilinxmultiregimpl145_regs0;
	builder_xilinxmultiregimpl146_regs0 <= main_inj_o_sys22;
	builder_xilinxmultiregimpl146_regs1 <= builder_xilinxmultiregimpl146_regs0;
	builder_xilinxmultiregimpl147_regs0 <= main_inj_o_sys23;
	builder_xilinxmultiregimpl147_regs1 <= builder_xilinxmultiregimpl147_regs0;
	builder_xilinxmultiregimpl148_regs0 <= main_inj_o_sys24;
	builder_xilinxmultiregimpl148_regs1 <= builder_xilinxmultiregimpl148_regs0;
	builder_xilinxmultiregimpl149_regs0 <= main_inj_o_sys25;
	builder_xilinxmultiregimpl149_regs1 <= builder_xilinxmultiregimpl149_regs0;
	builder_xilinxmultiregimpl150_regs0 <= main_inj_o_sys26;
	builder_xilinxmultiregimpl150_regs1 <= builder_xilinxmultiregimpl150_regs0;
	builder_xilinxmultiregimpl151_regs0 <= main_inj_o_sys27;
	builder_xilinxmultiregimpl151_regs1 <= builder_xilinxmultiregimpl151_regs0;
	builder_xilinxmultiregimpl152_regs0 <= main_inj_o_sys28;
	builder_xilinxmultiregimpl152_regs1 <= builder_xilinxmultiregimpl152_regs0;
	builder_xilinxmultiregimpl153_regs0 <= main_inj_o_sys29;
	builder_xilinxmultiregimpl153_regs1 <= builder_xilinxmultiregimpl153_regs0;
	builder_xilinxmultiregimpl154_regs0 <= main_inj_o_sys30;
	builder_xilinxmultiregimpl154_regs1 <= builder_xilinxmultiregimpl154_regs0;
	builder_xilinxmultiregimpl155_regs0 <= main_inj_o_sys31;
	builder_xilinxmultiregimpl155_regs1 <= builder_xilinxmultiregimpl155_regs0;
	builder_xilinxmultiregimpl156_regs0 <= main_inj_o_sys32;
	builder_xilinxmultiregimpl156_regs1 <= builder_xilinxmultiregimpl156_regs0;
	builder_xilinxmultiregimpl157_regs0 <= main_inj_o_sys33;
	builder_xilinxmultiregimpl157_regs1 <= builder_xilinxmultiregimpl157_regs0;
	builder_xilinxmultiregimpl158_regs0 <= main_inj_o_sys34;
	builder_xilinxmultiregimpl158_regs1 <= builder_xilinxmultiregimpl158_regs0;
	builder_xilinxmultiregimpl159_regs0 <= main_inj_o_sys35;
	builder_xilinxmultiregimpl159_regs1 <= builder_xilinxmultiregimpl159_regs0;
	builder_xilinxmultiregimpl160_regs0 <= main_inj_o_sys36;
	builder_xilinxmultiregimpl160_regs1 <= builder_xilinxmultiregimpl160_regs0;
	builder_xilinxmultiregimpl161_regs0 <= main_inj_o_sys37;
	builder_xilinxmultiregimpl161_regs1 <= builder_xilinxmultiregimpl161_regs0;
	builder_xilinxmultiregimpl162_regs0 <= main_inj_o_sys38;
	builder_xilinxmultiregimpl162_regs1 <= builder_xilinxmultiregimpl162_regs0;
	builder_xilinxmultiregimpl163_regs0 <= main_inj_o_sys39;
	builder_xilinxmultiregimpl163_regs1 <= builder_xilinxmultiregimpl163_regs0;
	builder_xilinxmultiregimpl164_regs0 <= main_inj_o_sys40;
	builder_xilinxmultiregimpl164_regs1 <= builder_xilinxmultiregimpl164_regs0;
	builder_xilinxmultiregimpl165_regs0 <= main_inj_o_sys41;
	builder_xilinxmultiregimpl165_regs1 <= builder_xilinxmultiregimpl165_regs0;
	builder_xilinxmultiregimpl166_regs0 <= main_inj_o_sys42;
	builder_xilinxmultiregimpl166_regs1 <= builder_xilinxmultiregimpl166_regs0;
	builder_xilinxmultiregimpl167_regs0 <= main_inj_o_sys43;
	builder_xilinxmultiregimpl167_regs1 <= builder_xilinxmultiregimpl167_regs0;
	builder_xilinxmultiregimpl168_regs0 <= main_inj_o_sys44;
	builder_xilinxmultiregimpl168_regs1 <= builder_xilinxmultiregimpl168_regs0;
	builder_xilinxmultiregimpl169_regs0 <= main_inj_o_sys45;
	builder_xilinxmultiregimpl169_regs1 <= builder_xilinxmultiregimpl169_regs0;
	builder_xilinxmultiregimpl170_regs0 <= main_inj_o_sys46;
	builder_xilinxmultiregimpl170_regs1 <= builder_xilinxmultiregimpl170_regs0;
	builder_xilinxmultiregimpl171_regs0 <= main_inj_o_sys47;
	builder_xilinxmultiregimpl171_regs1 <= builder_xilinxmultiregimpl171_regs0;
	builder_xilinxmultiregimpl172_regs0 <= main_inj_o_sys48;
	builder_xilinxmultiregimpl172_regs1 <= builder_xilinxmultiregimpl172_regs0;
	builder_xilinxmultiregimpl173_regs0 <= main_inj_o_sys49;
	builder_xilinxmultiregimpl173_regs1 <= builder_xilinxmultiregimpl173_regs0;
	builder_xilinxmultiregimpl174_regs0 <= main_inj_o_sys50;
	builder_xilinxmultiregimpl174_regs1 <= builder_xilinxmultiregimpl174_regs0;
	builder_xilinxmultiregimpl175_regs0 <= main_inj_o_sys51;
	builder_xilinxmultiregimpl175_regs1 <= builder_xilinxmultiregimpl175_regs0;
	builder_xilinxmultiregimpl176_regs0 <= main_inj_o_sys52;
	builder_xilinxmultiregimpl176_regs1 <= builder_xilinxmultiregimpl176_regs0;
	builder_xilinxmultiregimpl177_regs0 <= main_inj_o_sys53;
	builder_xilinxmultiregimpl177_regs1 <= builder_xilinxmultiregimpl177_regs0;
	builder_xilinxmultiregimpl178_regs0 <= main_inj_o_sys54;
	builder_xilinxmultiregimpl178_regs1 <= builder_xilinxmultiregimpl178_regs0;
	builder_xilinxmultiregimpl179_regs0 <= main_inj_o_sys55;
	builder_xilinxmultiregimpl179_regs1 <= builder_xilinxmultiregimpl179_regs0;
	builder_xilinxmultiregimpl180_regs0 <= main_inj_o_sys56;
	builder_xilinxmultiregimpl180_regs1 <= builder_xilinxmultiregimpl180_regs0;
	builder_xilinxmultiregimpl181_regs0 <= main_inj_o_sys57;
	builder_xilinxmultiregimpl181_regs1 <= builder_xilinxmultiregimpl181_regs0;
	builder_xilinxmultiregimpl182_regs0 <= main_inj_o_sys58;
	builder_xilinxmultiregimpl182_regs1 <= builder_xilinxmultiregimpl182_regs0;
	builder_xilinxmultiregimpl183_regs0 <= main_inj_o_sys59;
	builder_xilinxmultiregimpl183_regs1 <= builder_xilinxmultiregimpl183_regs0;
	builder_xilinxmultiregimpl184_regs0 <= main_inj_o_sys60;
	builder_xilinxmultiregimpl184_regs1 <= builder_xilinxmultiregimpl184_regs0;
	builder_xilinxmultiregimpl185_regs0 <= main_inj_o_sys61;
	builder_xilinxmultiregimpl185_regs1 <= builder_xilinxmultiregimpl185_regs0;
	builder_xilinxmultiregimpl186_regs0 <= main_inj_o_sys62;
	builder_xilinxmultiregimpl186_regs1 <= builder_xilinxmultiregimpl186_regs0;
	builder_xilinxmultiregimpl187_regs0 <= main_inj_o_sys63;
	builder_xilinxmultiregimpl187_regs1 <= builder_xilinxmultiregimpl187_regs0;
	builder_xilinxmultiregimpl188_regs0 <= main_inj_o_sys64;
	builder_xilinxmultiregimpl188_regs1 <= builder_xilinxmultiregimpl188_regs0;
	builder_xilinxmultiregimpl189_regs0 <= main_inj_o_sys65;
	builder_xilinxmultiregimpl189_regs1 <= builder_xilinxmultiregimpl189_regs0;
	builder_xilinxmultiregimpl190_regs0 <= main_inj_o_sys66;
	builder_xilinxmultiregimpl190_regs1 <= builder_xilinxmultiregimpl190_regs0;
	builder_xilinxmultiregimpl191_regs0 <= main_inj_o_sys67;
	builder_xilinxmultiregimpl191_regs1 <= builder_xilinxmultiregimpl191_regs0;
	builder_xilinxmultiregimpl192_regs0 <= main_inj_o_sys68;
	builder_xilinxmultiregimpl192_regs1 <= builder_xilinxmultiregimpl192_regs0;
	builder_xilinxmultiregimpl193_regs0 <= main_inj_o_sys69;
	builder_xilinxmultiregimpl193_regs1 <= builder_xilinxmultiregimpl193_regs0;
	builder_xilinxmultiregimpl194_regs0 <= main_inj_o_sys70;
	builder_xilinxmultiregimpl194_regs1 <= builder_xilinxmultiregimpl194_regs0;
	builder_xilinxmultiregimpl195_regs0 <= main_inj_o_sys71;
	builder_xilinxmultiregimpl195_regs1 <= builder_xilinxmultiregimpl195_regs0;
	builder_xilinxmultiregimpl196_regs0 <= main_inj_o_sys72;
	builder_xilinxmultiregimpl196_regs1 <= builder_xilinxmultiregimpl196_regs0;
	builder_xilinxmultiregimpl197_regs0 <= main_inj_o_sys73;
	builder_xilinxmultiregimpl197_regs1 <= builder_xilinxmultiregimpl197_regs0;
end

always @(posedge rio_phy_clk) begin
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd1))) begin
		main_inout_8x0_inout_8x0_oe_k <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_serdes_oe <= main_inout_8x0_inout_8x0_override_oe;
	end else begin
		main_inout_8x0_serdes_oe <= main_inout_8x0_inout_8x0_oe_k;
	end
	main_inout_8x0_inout_8x0_i_d <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_stb <= ((main_inout_8x0_inout_8x0_sample | (main_inout_8x0_inout_8x0_sensitivity[0] & (main_inout_8x0_serdes_i0[7] & (~main_inout_8x0_inout_8x0_i_d)))) | (main_inout_8x0_inout_8x0_sensitivity[1] & ((~main_inout_8x0_serdes_i0[7]) & main_inout_8x0_inout_8x0_i_d)));
	main_inout_8x0_inout_8x0_iinterface0_data <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_fine_ts <= main_inout_8x0_inout_8x0_o;
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0))) begin
		main_inout_8x0_inout_8x0_previous_data <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_override_o}};
	end else begin
		if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & (~main_inout_8x0_inout_8x0_previous_data)) & main_inout_8x0_inout_8x0_ointerface0_data[0])) begin
			main_inout_8x0_serdes_o0 <= builder_sync_f_t_array_muxed1;
		end else begin
			if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & main_inout_8x0_inout_8x0_previous_data) & (~main_inout_8x0_inout_8x0_ointerface0_data[0]))) begin
				main_inout_8x0_serdes_o0 <= builder_sync_f_t_array_muxed2;
			end else begin
				main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_previous_data}};
			end
		end
	end
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd1))) begin
		main_inout_8x1_inout_8x1_oe_k <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_serdes_oe <= main_inout_8x1_inout_8x1_override_oe;
	end else begin
		main_inout_8x1_serdes_oe <= main_inout_8x1_inout_8x1_oe_k;
	end
	main_inout_8x1_inout_8x1_i_d <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_stb <= ((main_inout_8x1_inout_8x1_sample | (main_inout_8x1_inout_8x1_sensitivity[0] & (main_inout_8x1_serdes_i0[7] & (~main_inout_8x1_inout_8x1_i_d)))) | (main_inout_8x1_inout_8x1_sensitivity[1] & ((~main_inout_8x1_serdes_i0[7]) & main_inout_8x1_inout_8x1_i_d)));
	main_inout_8x1_inout_8x1_iinterface1_data <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_fine_ts <= main_inout_8x1_inout_8x1_o;
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0))) begin
		main_inout_8x1_inout_8x1_previous_data <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_override_o}};
	end else begin
		if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & (~main_inout_8x1_inout_8x1_previous_data)) & main_inout_8x1_inout_8x1_ointerface1_data[0])) begin
			main_inout_8x1_serdes_o0 <= builder_sync_f_t_array_muxed3;
		end else begin
			if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & main_inout_8x1_inout_8x1_previous_data) & (~main_inout_8x1_inout_8x1_ointerface1_data[0]))) begin
				main_inout_8x1_serdes_o0 <= builder_sync_f_t_array_muxed4;
			end else begin
				main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_previous_data}};
			end
		end
	end
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd1))) begin
		main_inout_8x2_inout_8x2_oe_k <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_serdes_oe <= main_inout_8x2_inout_8x2_override_oe;
	end else begin
		main_inout_8x2_serdes_oe <= main_inout_8x2_inout_8x2_oe_k;
	end
	main_inout_8x2_inout_8x2_i_d <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_stb <= ((main_inout_8x2_inout_8x2_sample | (main_inout_8x2_inout_8x2_sensitivity[0] & (main_inout_8x2_serdes_i0[7] & (~main_inout_8x2_inout_8x2_i_d)))) | (main_inout_8x2_inout_8x2_sensitivity[1] & ((~main_inout_8x2_serdes_i0[7]) & main_inout_8x2_inout_8x2_i_d)));
	main_inout_8x2_inout_8x2_iinterface2_data <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_fine_ts <= main_inout_8x2_inout_8x2_o;
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0))) begin
		main_inout_8x2_inout_8x2_previous_data <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_override_o}};
	end else begin
		if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & (~main_inout_8x2_inout_8x2_previous_data)) & main_inout_8x2_inout_8x2_ointerface2_data[0])) begin
			main_inout_8x2_serdes_o0 <= builder_sync_f_t_array_muxed5;
		end else begin
			if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & main_inout_8x2_inout_8x2_previous_data) & (~main_inout_8x2_inout_8x2_ointerface2_data[0]))) begin
				main_inout_8x2_serdes_o0 <= builder_sync_f_t_array_muxed6;
			end else begin
				main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_previous_data}};
			end
		end
	end
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd1))) begin
		main_inout_8x3_inout_8x3_oe_k <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_serdes_oe <= main_inout_8x3_inout_8x3_override_oe;
	end else begin
		main_inout_8x3_serdes_oe <= main_inout_8x3_inout_8x3_oe_k;
	end
	main_inout_8x3_inout_8x3_i_d <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_stb <= ((main_inout_8x3_inout_8x3_sample | (main_inout_8x3_inout_8x3_sensitivity[0] & (main_inout_8x3_serdes_i0[7] & (~main_inout_8x3_inout_8x3_i_d)))) | (main_inout_8x3_inout_8x3_sensitivity[1] & ((~main_inout_8x3_serdes_i0[7]) & main_inout_8x3_inout_8x3_i_d)));
	main_inout_8x3_inout_8x3_iinterface3_data <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_fine_ts <= main_inout_8x3_inout_8x3_o;
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0))) begin
		main_inout_8x3_inout_8x3_previous_data <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_override_o}};
	end else begin
		if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & (~main_inout_8x3_inout_8x3_previous_data)) & main_inout_8x3_inout_8x3_ointerface3_data[0])) begin
			main_inout_8x3_serdes_o0 <= builder_sync_f_t_array_muxed7;
		end else begin
			if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & main_inout_8x3_inout_8x3_previous_data) & (~main_inout_8x3_inout_8x3_ointerface3_data[0]))) begin
				main_inout_8x3_serdes_o0 <= builder_sync_f_t_array_muxed8;
			end else begin
				main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_previous_data}};
			end
		end
	end
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd1))) begin
		main_inout_8x4_inout_8x4_oe_k <= main_inout_8x4_inout_8x4_ointerface4_data[0];
	end
	if (main_inout_8x4_inout_8x4_override_en) begin
		main_inout_8x4_serdes_oe <= main_inout_8x4_inout_8x4_override_oe;
	end else begin
		main_inout_8x4_serdes_oe <= main_inout_8x4_inout_8x4_oe_k;
	end
	main_inout_8x4_inout_8x4_i_d <= main_inout_8x4_serdes_i0[7];
	main_inout_8x4_inout_8x4_iinterface4_stb <= ((main_inout_8x4_inout_8x4_sample | (main_inout_8x4_inout_8x4_sensitivity[0] & (main_inout_8x4_serdes_i0[7] & (~main_inout_8x4_inout_8x4_i_d)))) | (main_inout_8x4_inout_8x4_sensitivity[1] & ((~main_inout_8x4_serdes_i0[7]) & main_inout_8x4_inout_8x4_i_d)));
	main_inout_8x4_inout_8x4_iinterface4_data <= main_inout_8x4_serdes_i0[7];
	main_inout_8x4_inout_8x4_iinterface4_fine_ts <= main_inout_8x4_inout_8x4_o;
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0))) begin
		main_inout_8x4_inout_8x4_previous_data <= main_inout_8x4_inout_8x4_ointerface4_data[0];
	end
	if (main_inout_8x4_inout_8x4_override_en) begin
		main_inout_8x4_serdes_o0 <= {8{main_inout_8x4_inout_8x4_override_o}};
	end else begin
		if ((((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0)) & (~main_inout_8x4_inout_8x4_previous_data)) & main_inout_8x4_inout_8x4_ointerface4_data[0])) begin
			main_inout_8x4_serdes_o0 <= builder_sync_f_t_array_muxed9;
		end else begin
			if ((((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0)) & main_inout_8x4_inout_8x4_previous_data) & (~main_inout_8x4_inout_8x4_ointerface4_data[0]))) begin
				main_inout_8x4_serdes_o0 <= builder_sync_f_t_array_muxed10;
			end else begin
				main_inout_8x4_serdes_o0 <= {8{main_inout_8x4_inout_8x4_previous_data}};
			end
		end
	end
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd1))) begin
		main_inout_8x5_inout_8x5_oe_k <= main_inout_8x5_inout_8x5_ointerface5_data[0];
	end
	if (main_inout_8x5_inout_8x5_override_en) begin
		main_inout_8x5_serdes_oe <= main_inout_8x5_inout_8x5_override_oe;
	end else begin
		main_inout_8x5_serdes_oe <= main_inout_8x5_inout_8x5_oe_k;
	end
	main_inout_8x5_inout_8x5_i_d <= main_inout_8x5_serdes_i0[7];
	main_inout_8x5_inout_8x5_iinterface5_stb <= ((main_inout_8x5_inout_8x5_sample | (main_inout_8x5_inout_8x5_sensitivity[0] & (main_inout_8x5_serdes_i0[7] & (~main_inout_8x5_inout_8x5_i_d)))) | (main_inout_8x5_inout_8x5_sensitivity[1] & ((~main_inout_8x5_serdes_i0[7]) & main_inout_8x5_inout_8x5_i_d)));
	main_inout_8x5_inout_8x5_iinterface5_data <= main_inout_8x5_serdes_i0[7];
	main_inout_8x5_inout_8x5_iinterface5_fine_ts <= main_inout_8x5_inout_8x5_o;
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0))) begin
		main_inout_8x5_inout_8x5_previous_data <= main_inout_8x5_inout_8x5_ointerface5_data[0];
	end
	if (main_inout_8x5_inout_8x5_override_en) begin
		main_inout_8x5_serdes_o0 <= {8{main_inout_8x5_inout_8x5_override_o}};
	end else begin
		if ((((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0)) & (~main_inout_8x5_inout_8x5_previous_data)) & main_inout_8x5_inout_8x5_ointerface5_data[0])) begin
			main_inout_8x5_serdes_o0 <= builder_sync_f_t_array_muxed11;
		end else begin
			if ((((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0)) & main_inout_8x5_inout_8x5_previous_data) & (~main_inout_8x5_inout_8x5_ointerface5_data[0]))) begin
				main_inout_8x5_serdes_o0 <= builder_sync_f_t_array_muxed12;
			end else begin
				main_inout_8x5_serdes_o0 <= {8{main_inout_8x5_inout_8x5_previous_data}};
			end
		end
	end
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd1))) begin
		main_inout_8x6_inout_8x6_oe_k <= main_inout_8x6_inout_8x6_ointerface6_data[0];
	end
	if (main_inout_8x6_inout_8x6_override_en) begin
		main_inout_8x6_serdes_oe <= main_inout_8x6_inout_8x6_override_oe;
	end else begin
		main_inout_8x6_serdes_oe <= main_inout_8x6_inout_8x6_oe_k;
	end
	main_inout_8x6_inout_8x6_i_d <= main_inout_8x6_serdes_i0[7];
	main_inout_8x6_inout_8x6_iinterface6_stb <= ((main_inout_8x6_inout_8x6_sample | (main_inout_8x6_inout_8x6_sensitivity[0] & (main_inout_8x6_serdes_i0[7] & (~main_inout_8x6_inout_8x6_i_d)))) | (main_inout_8x6_inout_8x6_sensitivity[1] & ((~main_inout_8x6_serdes_i0[7]) & main_inout_8x6_inout_8x6_i_d)));
	main_inout_8x6_inout_8x6_iinterface6_data <= main_inout_8x6_serdes_i0[7];
	main_inout_8x6_inout_8x6_iinterface6_fine_ts <= main_inout_8x6_inout_8x6_o;
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0))) begin
		main_inout_8x6_inout_8x6_previous_data <= main_inout_8x6_inout_8x6_ointerface6_data[0];
	end
	if (main_inout_8x6_inout_8x6_override_en) begin
		main_inout_8x6_serdes_o0 <= {8{main_inout_8x6_inout_8x6_override_o}};
	end else begin
		if ((((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0)) & (~main_inout_8x6_inout_8x6_previous_data)) & main_inout_8x6_inout_8x6_ointerface6_data[0])) begin
			main_inout_8x6_serdes_o0 <= builder_sync_f_t_array_muxed13;
		end else begin
			if ((((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0)) & main_inout_8x6_inout_8x6_previous_data) & (~main_inout_8x6_inout_8x6_ointerface6_data[0]))) begin
				main_inout_8x6_serdes_o0 <= builder_sync_f_t_array_muxed14;
			end else begin
				main_inout_8x6_serdes_o0 <= {8{main_inout_8x6_inout_8x6_previous_data}};
			end
		end
	end
	if ((main_inout_8x7_inout_8x7_ointerface7_stb & (main_inout_8x7_inout_8x7_ointerface7_address == 1'd1))) begin
		main_inout_8x7_inout_8x7_oe_k <= main_inout_8x7_inout_8x7_ointerface7_data[0];
	end
	if (main_inout_8x7_inout_8x7_override_en) begin
		main_inout_8x7_serdes_oe <= main_inout_8x7_inout_8x7_override_oe;
	end else begin
		main_inout_8x7_serdes_oe <= main_inout_8x7_inout_8x7_oe_k;
	end
	main_inout_8x7_inout_8x7_i_d <= main_inout_8x7_serdes_i0[7];
	main_inout_8x7_inout_8x7_iinterface7_stb <= ((main_inout_8x7_inout_8x7_sample | (main_inout_8x7_inout_8x7_sensitivity[0] & (main_inout_8x7_serdes_i0[7] & (~main_inout_8x7_inout_8x7_i_d)))) | (main_inout_8x7_inout_8x7_sensitivity[1] & ((~main_inout_8x7_serdes_i0[7]) & main_inout_8x7_inout_8x7_i_d)));
	main_inout_8x7_inout_8x7_iinterface7_data <= main_inout_8x7_serdes_i0[7];
	main_inout_8x7_inout_8x7_iinterface7_fine_ts <= main_inout_8x7_inout_8x7_o;
	if ((main_inout_8x7_inout_8x7_ointerface7_stb & (main_inout_8x7_inout_8x7_ointerface7_address == 1'd0))) begin
		main_inout_8x7_inout_8x7_previous_data <= main_inout_8x7_inout_8x7_ointerface7_data[0];
	end
	if (main_inout_8x7_inout_8x7_override_en) begin
		main_inout_8x7_serdes_o0 <= {8{main_inout_8x7_inout_8x7_override_o}};
	end else begin
		if ((((main_inout_8x7_inout_8x7_ointerface7_stb & (main_inout_8x7_inout_8x7_ointerface7_address == 1'd0)) & (~main_inout_8x7_inout_8x7_previous_data)) & main_inout_8x7_inout_8x7_ointerface7_data[0])) begin
			main_inout_8x7_serdes_o0 <= builder_sync_f_t_array_muxed15;
		end else begin
			if ((((main_inout_8x7_inout_8x7_ointerface7_stb & (main_inout_8x7_inout_8x7_ointerface7_address == 1'd0)) & main_inout_8x7_inout_8x7_previous_data) & (~main_inout_8x7_inout_8x7_ointerface7_data[0]))) begin
				main_inout_8x7_serdes_o0 <= builder_sync_f_t_array_muxed16;
			end else begin
				main_inout_8x7_serdes_o0 <= {8{main_inout_8x7_inout_8x7_previous_data}};
			end
		end
	end
	if (main_output_8x0_stb) begin
		main_output_8x0_previous_data <= main_output_8x0_data;
	end
	if (main_output_8x0_override_en) begin
		main_output_8x0_o <= {8{main_output_8x0_override_o}};
	end else begin
		if (((main_output_8x0_stb & (~main_output_8x0_previous_data)) & main_output_8x0_data)) begin
			main_output_8x0_o <= builder_sync_f_t_array_muxed17;
		end else begin
			if (((main_output_8x0_stb & main_output_8x0_previous_data) & (~main_output_8x0_data))) begin
				main_output_8x0_o <= builder_sync_f_t_array_muxed18;
			end else begin
				main_output_8x0_o <= {8{main_output_8x0_previous_data}};
			end
		end
	end
	if (main_output_8x1_stb) begin
		main_output_8x1_previous_data <= main_output_8x1_data;
	end
	if (main_output_8x1_override_en) begin
		main_output_8x1_o <= {8{main_output_8x1_override_o}};
	end else begin
		if (((main_output_8x1_stb & (~main_output_8x1_previous_data)) & main_output_8x1_data)) begin
			main_output_8x1_o <= builder_sync_f_t_array_muxed19;
		end else begin
			if (((main_output_8x1_stb & main_output_8x1_previous_data) & (~main_output_8x1_data))) begin
				main_output_8x1_o <= builder_sync_f_t_array_muxed20;
			end else begin
				main_output_8x1_o <= {8{main_output_8x1_previous_data}};
			end
		end
	end
	if (main_output_8x2_stb) begin
		main_output_8x2_previous_data <= main_output_8x2_data;
	end
	if (main_output_8x2_override_en) begin
		main_output_8x2_o <= {8{main_output_8x2_override_o}};
	end else begin
		if (((main_output_8x2_stb & (~main_output_8x2_previous_data)) & main_output_8x2_data)) begin
			main_output_8x2_o <= builder_sync_f_t_array_muxed21;
		end else begin
			if (((main_output_8x2_stb & main_output_8x2_previous_data) & (~main_output_8x2_data))) begin
				main_output_8x2_o <= builder_sync_f_t_array_muxed22;
			end else begin
				main_output_8x2_o <= {8{main_output_8x2_previous_data}};
			end
		end
	end
	if (main_output_8x3_stb) begin
		main_output_8x3_previous_data <= main_output_8x3_data;
	end
	if (main_output_8x3_override_en) begin
		main_output_8x3_o <= {8{main_output_8x3_override_o}};
	end else begin
		if (((main_output_8x3_stb & (~main_output_8x3_previous_data)) & main_output_8x3_data)) begin
			main_output_8x3_o <= builder_sync_f_t_array_muxed23;
		end else begin
			if (((main_output_8x3_stb & main_output_8x3_previous_data) & (~main_output_8x3_data))) begin
				main_output_8x3_o <= builder_sync_f_t_array_muxed24;
			end else begin
				main_output_8x3_o <= {8{main_output_8x3_previous_data}};
			end
		end
	end
	if (main_output_8x4_stb) begin
		main_output_8x4_previous_data <= main_output_8x4_data;
	end
	if (main_output_8x4_override_en) begin
		main_output_8x4_o <= {8{main_output_8x4_override_o}};
	end else begin
		if (((main_output_8x4_stb & (~main_output_8x4_previous_data)) & main_output_8x4_data)) begin
			main_output_8x4_o <= builder_sync_f_t_array_muxed25;
		end else begin
			if (((main_output_8x4_stb & main_output_8x4_previous_data) & (~main_output_8x4_data))) begin
				main_output_8x4_o <= builder_sync_f_t_array_muxed26;
			end else begin
				main_output_8x4_o <= {8{main_output_8x4_previous_data}};
			end
		end
	end
	if (main_output_8x5_stb) begin
		main_output_8x5_previous_data <= main_output_8x5_data;
	end
	if (main_output_8x5_override_en) begin
		main_output_8x5_o <= {8{main_output_8x5_override_o}};
	end else begin
		if (((main_output_8x5_stb & (~main_output_8x5_previous_data)) & main_output_8x5_data)) begin
			main_output_8x5_o <= builder_sync_f_t_array_muxed27;
		end else begin
			if (((main_output_8x5_stb & main_output_8x5_previous_data) & (~main_output_8x5_data))) begin
				main_output_8x5_o <= builder_sync_f_t_array_muxed28;
			end else begin
				main_output_8x5_o <= {8{main_output_8x5_previous_data}};
			end
		end
	end
	if (main_output_8x6_stb) begin
		main_output_8x6_previous_data <= main_output_8x6_data;
	end
	if (main_output_8x6_override_en) begin
		main_output_8x6_o <= {8{main_output_8x6_override_o}};
	end else begin
		if (((main_output_8x6_stb & (~main_output_8x6_previous_data)) & main_output_8x6_data)) begin
			main_output_8x6_o <= builder_sync_f_t_array_muxed29;
		end else begin
			if (((main_output_8x6_stb & main_output_8x6_previous_data) & (~main_output_8x6_data))) begin
				main_output_8x6_o <= builder_sync_f_t_array_muxed30;
			end else begin
				main_output_8x6_o <= {8{main_output_8x6_previous_data}};
			end
		end
	end
	if (main_output_8x7_stb) begin
		main_output_8x7_previous_data <= main_output_8x7_data;
	end
	if (main_output_8x7_override_en) begin
		main_output_8x7_o <= {8{main_output_8x7_override_o}};
	end else begin
		if (((main_output_8x7_stb & (~main_output_8x7_previous_data)) & main_output_8x7_data)) begin
			main_output_8x7_o <= builder_sync_f_t_array_muxed31;
		end else begin
			if (((main_output_8x7_stb & main_output_8x7_previous_data) & (~main_output_8x7_data))) begin
				main_output_8x7_o <= builder_sync_f_t_array_muxed32;
			end else begin
				main_output_8x7_o <= {8{main_output_8x7_previous_data}};
			end
		end
	end
	if (main_spimaster0_iinterface0_stb) begin
		main_spimaster0_read <= 1'd0;
	end
	if ((main_spimaster0_ointerface0_stb & main_spimaster0_spimachine0_writable)) begin
		if (main_spimaster0_ointerface0_address) begin
			{main_spimaster0_config_cs, main_spimaster0_config_div, main_spimaster0_config_padding, main_spimaster0_config_length, main_spimaster0_config_half_duplex, main_spimaster0_config_lsb_first, main_spimaster0_config_clk_phase, main_spimaster0_config_clk_polarity, main_spimaster0_config_cs_polarity, main_spimaster0_config_input, main_spimaster0_config_end, main_spimaster0_config_offline} <= main_spimaster0_ointerface0_data;
		end else begin
			main_spimaster0_read <= main_spimaster0_config_input;
		end
	end
	if (main_spimaster0_interface_ce) begin
		main_spimaster0_interface_cs1 <= (({3{main_spimaster0_interface_cs_next}} & main_spimaster0_interface_cs0) ^ (~main_spimaster0_interface_cs_polarity));
		main_spimaster0_interface_clk <= (main_spimaster0_interface_clk_next ^ main_spimaster0_interface_clk_polarity);
	end
	if (main_spimaster0_interface_sample) begin
		main_spimaster0_interface_miso_reg <= main_spimaster0_interface_miso;
		main_spimaster0_interface_mosi_reg <= main_spimaster0_interface_mosi;
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_n <= main_spimaster0_spimachine0_length;
		main_spimaster0_spimachine0_end1 <= main_spimaster0_spimachine0_end0;
	end
	if (main_spimaster0_spimachine0_shift) begin
		main_spimaster0_spimachine0_n <= (main_spimaster0_spimachine0_n - 1'd1);
	end
	if (main_spimaster0_spimachine0_shift) begin
		main_spimaster0_spimachine0_sr <= main_spimaster0_spimachine0_pdi;
		main_spimaster0_spimachine0_sdo <= (main_spimaster0_spimachine0_lsb_first ? main_spimaster0_spimachine0_pdi[0] : main_spimaster0_spimachine0_pdi[31]);
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_sr <= main_spimaster0_spimachine0_pdo;
		main_spimaster0_spimachine0_sdo <= (main_spimaster0_spimachine0_lsb_first ? main_spimaster0_spimachine0_pdo[0] : main_spimaster0_spimachine0_pdo[31]);
	end
	if (main_spimaster0_spimachine0_count) begin
		if (main_spimaster0_spimachine0_cnt_done) begin
			if (main_spimaster0_spimachine0_do_extend) begin
				main_spimaster0_spimachine0_do_extend <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_cnt <= main_spimaster0_spimachine0_div[7:1];
				main_spimaster0_spimachine0_do_extend <= (main_spimaster0_spimachine0_extend & main_spimaster0_spimachine0_div[0]);
			end
		end else begin
			main_spimaster0_spimachine0_cnt <= (main_spimaster0_spimachine0_cnt - 1'd1);
		end
	end
	builder_spimaster0_state <= builder_spimaster0_next_state;
	if (main_output_8x8_stb) begin
		main_output_8x8_previous_data <= main_output_8x8_data;
	end
	if (main_output_8x8_override_en) begin
		main_output_8x8_o <= {8{main_output_8x8_override_o}};
	end else begin
		if (((main_output_8x8_stb & (~main_output_8x8_previous_data)) & main_output_8x8_data)) begin
			main_output_8x8_o <= builder_sync_f_t_array_muxed33;
		end else begin
			if (((main_output_8x8_stb & main_output_8x8_previous_data) & (~main_output_8x8_data))) begin
				main_output_8x8_o <= builder_sync_f_t_array_muxed34;
			end else begin
				main_output_8x8_o <= {8{main_output_8x8_previous_data}};
			end
		end
	end
	if (main_output_8x9_stb) begin
		main_output_8x9_previous_data <= main_output_8x9_data;
	end
	if (main_output_8x9_override_en) begin
		main_output_8x9_o <= {8{main_output_8x9_override_o}};
	end else begin
		if (((main_output_8x9_stb & (~main_output_8x9_previous_data)) & main_output_8x9_data)) begin
			main_output_8x9_o <= builder_sync_f_t_array_muxed35;
		end else begin
			if (((main_output_8x9_stb & main_output_8x9_previous_data) & (~main_output_8x9_data))) begin
				main_output_8x9_o <= builder_sync_f_t_array_muxed36;
			end else begin
				main_output_8x9_o <= {8{main_output_8x9_previous_data}};
			end
		end
	end
	if (main_output_8x10_stb) begin
		main_output_8x10_previous_data <= main_output_8x10_data;
	end
	if (main_output_8x10_override_en) begin
		main_output_8x10_o <= {8{main_output_8x10_override_o}};
	end else begin
		if (((main_output_8x10_stb & (~main_output_8x10_previous_data)) & main_output_8x10_data)) begin
			main_output_8x10_o <= builder_sync_f_t_array_muxed37;
		end else begin
			if (((main_output_8x10_stb & main_output_8x10_previous_data) & (~main_output_8x10_data))) begin
				main_output_8x10_o <= builder_sync_f_t_array_muxed38;
			end else begin
				main_output_8x10_o <= {8{main_output_8x10_previous_data}};
			end
		end
	end
	if (main_output_8x11_stb) begin
		main_output_8x11_previous_data <= main_output_8x11_data;
	end
	if (main_output_8x11_override_en) begin
		main_output_8x11_o <= {8{main_output_8x11_override_o}};
	end else begin
		if (((main_output_8x11_stb & (~main_output_8x11_previous_data)) & main_output_8x11_data)) begin
			main_output_8x11_o <= builder_sync_f_t_array_muxed39;
		end else begin
			if (((main_output_8x11_stb & main_output_8x11_previous_data) & (~main_output_8x11_data))) begin
				main_output_8x11_o <= builder_sync_f_t_array_muxed40;
			end else begin
				main_output_8x11_o <= {8{main_output_8x11_previous_data}};
			end
		end
	end
	if (main_output_8x12_stb) begin
		main_output_8x12_previous_data <= main_output_8x12_data;
	end
	if (main_output_8x12_override_en) begin
		main_output_8x12_o <= {8{main_output_8x12_override_o}};
	end else begin
		if (((main_output_8x12_stb & (~main_output_8x12_previous_data)) & main_output_8x12_data)) begin
			main_output_8x12_o <= builder_sync_f_t_array_muxed41;
		end else begin
			if (((main_output_8x12_stb & main_output_8x12_previous_data) & (~main_output_8x12_data))) begin
				main_output_8x12_o <= builder_sync_f_t_array_muxed42;
			end else begin
				main_output_8x12_o <= {8{main_output_8x12_previous_data}};
			end
		end
	end
	if (main_spimaster1_iinterface1_stb) begin
		main_spimaster1_read <= 1'd0;
	end
	if ((main_spimaster1_ointerface1_stb & main_spimaster1_spimachine1_writable)) begin
		if (main_spimaster1_ointerface1_address) begin
			{main_spimaster1_config_cs, main_spimaster1_config_div, main_spimaster1_config_padding, main_spimaster1_config_length, main_spimaster1_config_half_duplex, main_spimaster1_config_lsb_first, main_spimaster1_config_clk_phase, main_spimaster1_config_clk_polarity, main_spimaster1_config_cs_polarity, main_spimaster1_config_input, main_spimaster1_config_end, main_spimaster1_config_offline} <= main_spimaster1_ointerface1_data;
		end else begin
			main_spimaster1_read <= main_spimaster1_config_input;
		end
	end
	if (main_spimaster1_interface_ce) begin
		main_spimaster1_interface_cs1 <= (({3{main_spimaster1_interface_cs_next}} & main_spimaster1_interface_cs0) ^ (~main_spimaster1_interface_cs_polarity));
		main_spimaster1_interface_clk <= (main_spimaster1_interface_clk_next ^ main_spimaster1_interface_clk_polarity);
	end
	if (main_spimaster1_interface_sample) begin
		main_spimaster1_interface_miso_reg <= main_spimaster1_interface_miso;
		main_spimaster1_interface_mosi_reg <= main_spimaster1_interface_mosi;
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_n <= main_spimaster1_spimachine1_length;
		main_spimaster1_spimachine1_end1 <= main_spimaster1_spimachine1_end0;
	end
	if (main_spimaster1_spimachine1_shift) begin
		main_spimaster1_spimachine1_n <= (main_spimaster1_spimachine1_n - 1'd1);
	end
	if (main_spimaster1_spimachine1_shift) begin
		main_spimaster1_spimachine1_sr <= main_spimaster1_spimachine1_pdi;
		main_spimaster1_spimachine1_sdo <= (main_spimaster1_spimachine1_lsb_first ? main_spimaster1_spimachine1_pdi[0] : main_spimaster1_spimachine1_pdi[31]);
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_sr <= main_spimaster1_spimachine1_pdo;
		main_spimaster1_spimachine1_sdo <= (main_spimaster1_spimachine1_lsb_first ? main_spimaster1_spimachine1_pdo[0] : main_spimaster1_spimachine1_pdo[31]);
	end
	if (main_spimaster1_spimachine1_count) begin
		if (main_spimaster1_spimachine1_cnt_done) begin
			if (main_spimaster1_spimachine1_do_extend) begin
				main_spimaster1_spimachine1_do_extend <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_cnt <= main_spimaster1_spimachine1_div[7:1];
				main_spimaster1_spimachine1_do_extend <= (main_spimaster1_spimachine1_extend & main_spimaster1_spimachine1_div[0]);
			end
		end else begin
			main_spimaster1_spimachine1_cnt <= (main_spimaster1_spimachine1_cnt - 1'd1);
		end
	end
	builder_spimaster1_state <= builder_spimaster1_next_state;
	if (main_output_8x13_stb) begin
		main_output_8x13_previous_data <= main_output_8x13_data;
	end
	if (main_output_8x13_override_en) begin
		main_output_8x13_o <= {8{main_output_8x13_override_o}};
	end else begin
		if (((main_output_8x13_stb & (~main_output_8x13_previous_data)) & main_output_8x13_data)) begin
			main_output_8x13_o <= builder_sync_f_t_array_muxed43;
		end else begin
			if (((main_output_8x13_stb & main_output_8x13_previous_data) & (~main_output_8x13_data))) begin
				main_output_8x13_o <= builder_sync_f_t_array_muxed44;
			end else begin
				main_output_8x13_o <= {8{main_output_8x13_previous_data}};
			end
		end
	end
	if (main_output_8x14_stb) begin
		main_output_8x14_previous_data <= main_output_8x14_data;
	end
	if (main_output_8x14_override_en) begin
		main_output_8x14_o <= {8{main_output_8x14_override_o}};
	end else begin
		if (((main_output_8x14_stb & (~main_output_8x14_previous_data)) & main_output_8x14_data)) begin
			main_output_8x14_o <= builder_sync_f_t_array_muxed45;
		end else begin
			if (((main_output_8x14_stb & main_output_8x14_previous_data) & (~main_output_8x14_data))) begin
				main_output_8x14_o <= builder_sync_f_t_array_muxed46;
			end else begin
				main_output_8x14_o <= {8{main_output_8x14_previous_data}};
			end
		end
	end
	if (main_output_8x15_stb) begin
		main_output_8x15_previous_data <= main_output_8x15_data;
	end
	if (main_output_8x15_override_en) begin
		main_output_8x15_o <= {8{main_output_8x15_override_o}};
	end else begin
		if (((main_output_8x15_stb & (~main_output_8x15_previous_data)) & main_output_8x15_data)) begin
			main_output_8x15_o <= builder_sync_f_t_array_muxed47;
		end else begin
			if (((main_output_8x15_stb & main_output_8x15_previous_data) & (~main_output_8x15_data))) begin
				main_output_8x15_o <= builder_sync_f_t_array_muxed48;
			end else begin
				main_output_8x15_o <= {8{main_output_8x15_previous_data}};
			end
		end
	end
	if (main_output_8x16_stb) begin
		main_output_8x16_previous_data <= main_output_8x16_data;
	end
	if (main_output_8x16_override_en) begin
		main_output_8x16_o <= {8{main_output_8x16_override_o}};
	end else begin
		if (((main_output_8x16_stb & (~main_output_8x16_previous_data)) & main_output_8x16_data)) begin
			main_output_8x16_o <= builder_sync_f_t_array_muxed49;
		end else begin
			if (((main_output_8x16_stb & main_output_8x16_previous_data) & (~main_output_8x16_data))) begin
				main_output_8x16_o <= builder_sync_f_t_array_muxed50;
			end else begin
				main_output_8x16_o <= {8{main_output_8x16_previous_data}};
			end
		end
	end
	if (main_output_8x17_stb) begin
		main_output_8x17_previous_data <= main_output_8x17_data;
	end
	if (main_output_8x17_override_en) begin
		main_output_8x17_o <= {8{main_output_8x17_override_o}};
	end else begin
		if (((main_output_8x17_stb & (~main_output_8x17_previous_data)) & main_output_8x17_data)) begin
			main_output_8x17_o <= builder_sync_f_t_array_muxed51;
		end else begin
			if (((main_output_8x17_stb & main_output_8x17_previous_data) & (~main_output_8x17_data))) begin
				main_output_8x17_o <= builder_sync_f_t_array_muxed52;
			end else begin
				main_output_8x17_o <= {8{main_output_8x17_previous_data}};
			end
		end
	end
	if (main_spimaster2_iinterface2_stb) begin
		main_spimaster2_read <= 1'd0;
	end
	if ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable)) begin
		if (main_spimaster2_ointerface2_address) begin
			{main_spimaster2_config_cs, main_spimaster2_config_div, main_spimaster2_config_padding, main_spimaster2_config_length, main_spimaster2_config_half_duplex, main_spimaster2_config_lsb_first, main_spimaster2_config_clk_phase, main_spimaster2_config_clk_polarity, main_spimaster2_config_cs_polarity, main_spimaster2_config_input, main_spimaster2_config_end, main_spimaster2_config_offline} <= main_spimaster2_ointerface2_data;
		end else begin
			main_spimaster2_read <= main_spimaster2_config_input;
		end
	end
	if (main_spimaster2_interface_ce) begin
		main_spimaster2_interface_cs1 <= (({3{main_spimaster2_interface_cs_next}} & main_spimaster2_interface_cs0) ^ (~main_spimaster2_interface_cs_polarity));
		main_spimaster2_interface_clk <= (main_spimaster2_interface_clk_next ^ main_spimaster2_interface_clk_polarity);
	end
	if (main_spimaster2_interface_sample) begin
		main_spimaster2_interface_miso_reg <= main_spimaster2_interface_miso;
		main_spimaster2_interface_mosi_reg <= main_spimaster2_interface_mosi;
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_n <= main_spimaster2_spimachine2_length;
		main_spimaster2_spimachine2_end1 <= main_spimaster2_spimachine2_end0;
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_n <= (main_spimaster2_spimachine2_n - 1'd1);
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdi;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdi[0] : main_spimaster2_spimachine2_pdi[31]);
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdo;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdo[0] : main_spimaster2_spimachine2_pdo[31]);
	end
	if (main_spimaster2_spimachine2_count) begin
		if (main_spimaster2_spimachine2_cnt_done) begin
			if (main_spimaster2_spimachine2_do_extend) begin
				main_spimaster2_spimachine2_do_extend <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_cnt <= main_spimaster2_spimachine2_div[7:1];
				main_spimaster2_spimachine2_do_extend <= (main_spimaster2_spimachine2_extend & main_spimaster2_spimachine2_div[0]);
			end
		end else begin
			main_spimaster2_spimachine2_cnt <= (main_spimaster2_spimachine2_cnt - 1'd1);
		end
	end
	builder_spimaster2_state <= builder_spimaster2_next_state;
	if (main_output_8x18_stb) begin
		main_output_8x18_previous_data <= main_output_8x18_data;
	end
	if (main_output_8x18_override_en) begin
		main_output_8x18_o <= {8{main_output_8x18_override_o}};
	end else begin
		if (((main_output_8x18_stb & (~main_output_8x18_previous_data)) & main_output_8x18_data)) begin
			main_output_8x18_o <= builder_sync_f_t_array_muxed53;
		end else begin
			if (((main_output_8x18_stb & main_output_8x18_previous_data) & (~main_output_8x18_data))) begin
				main_output_8x18_o <= builder_sync_f_t_array_muxed54;
			end else begin
				main_output_8x18_o <= {8{main_output_8x18_previous_data}};
			end
		end
	end
	if (main_output_8x19_stb) begin
		main_output_8x19_previous_data <= main_output_8x19_data;
	end
	if (main_output_8x19_override_en) begin
		main_output_8x19_o <= {8{main_output_8x19_override_o}};
	end else begin
		if (((main_output_8x19_stb & (~main_output_8x19_previous_data)) & main_output_8x19_data)) begin
			main_output_8x19_o <= builder_sync_f_t_array_muxed55;
		end else begin
			if (((main_output_8x19_stb & main_output_8x19_previous_data) & (~main_output_8x19_data))) begin
				main_output_8x19_o <= builder_sync_f_t_array_muxed56;
			end else begin
				main_output_8x19_o <= {8{main_output_8x19_previous_data}};
			end
		end
	end
	if (main_output_8x20_stb) begin
		main_output_8x20_previous_data <= main_output_8x20_data;
	end
	if (main_output_8x20_override_en) begin
		main_output_8x20_o <= {8{main_output_8x20_override_o}};
	end else begin
		if (((main_output_8x20_stb & (~main_output_8x20_previous_data)) & main_output_8x20_data)) begin
			main_output_8x20_o <= builder_sync_f_t_array_muxed57;
		end else begin
			if (((main_output_8x20_stb & main_output_8x20_previous_data) & (~main_output_8x20_data))) begin
				main_output_8x20_o <= builder_sync_f_t_array_muxed58;
			end else begin
				main_output_8x20_o <= {8{main_output_8x20_previous_data}};
			end
		end
	end
	if (main_output_8x21_stb) begin
		main_output_8x21_previous_data <= main_output_8x21_data;
	end
	if (main_output_8x21_override_en) begin
		main_output_8x21_o <= {8{main_output_8x21_override_o}};
	end else begin
		if (((main_output_8x21_stb & (~main_output_8x21_previous_data)) & main_output_8x21_data)) begin
			main_output_8x21_o <= builder_sync_f_t_array_muxed59;
		end else begin
			if (((main_output_8x21_stb & main_output_8x21_previous_data) & (~main_output_8x21_data))) begin
				main_output_8x21_o <= builder_sync_f_t_array_muxed60;
			end else begin
				main_output_8x21_o <= {8{main_output_8x21_previous_data}};
			end
		end
	end
	if (main_output_8x22_stb) begin
		main_output_8x22_previous_data <= main_output_8x22_data;
	end
	if (main_output_8x22_override_en) begin
		main_output_8x22_o <= {8{main_output_8x22_override_o}};
	end else begin
		if (((main_output_8x22_stb & (~main_output_8x22_previous_data)) & main_output_8x22_data)) begin
			main_output_8x22_o <= builder_sync_f_t_array_muxed61;
		end else begin
			if (((main_output_8x22_stb & main_output_8x22_previous_data) & (~main_output_8x22_data))) begin
				main_output_8x22_o <= builder_sync_f_t_array_muxed62;
			end else begin
				main_output_8x22_o <= {8{main_output_8x22_previous_data}};
			end
		end
	end
	if (main_output0_stb) begin
		main_output0_pad_k <= main_output0_data;
	end
	if (main_output0_override_en) begin
		main_output0_pad_o <= main_output0_override_o;
	end else begin
		main_output0_pad_o <= main_output0_pad_k;
	end
	if (main_output1_stb) begin
		main_output1_pad_k <= main_output1_data;
	end
	if (main_output1_override_en) begin
		main_output1_pad_o <= main_output1_override_o;
	end else begin
		main_output1_pad_o <= main_output1_pad_k;
	end
	if (rio_phy_rst) begin
		main_inout_8x0_serdes_o0 <= 8'd0;
		main_inout_8x0_serdes_oe <= 1'd0;
		main_inout_8x0_inout_8x0_iinterface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_previous_data <= 1'd0;
		main_inout_8x0_inout_8x0_oe_k <= 1'd0;
		main_inout_8x0_inout_8x0_i_d <= 1'd0;
		main_inout_8x1_serdes_o0 <= 8'd0;
		main_inout_8x1_serdes_oe <= 1'd0;
		main_inout_8x1_inout_8x1_iinterface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_previous_data <= 1'd0;
		main_inout_8x1_inout_8x1_oe_k <= 1'd0;
		main_inout_8x1_inout_8x1_i_d <= 1'd0;
		main_inout_8x2_serdes_o0 <= 8'd0;
		main_inout_8x2_serdes_oe <= 1'd0;
		main_inout_8x2_inout_8x2_iinterface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_previous_data <= 1'd0;
		main_inout_8x2_inout_8x2_oe_k <= 1'd0;
		main_inout_8x2_inout_8x2_i_d <= 1'd0;
		main_inout_8x3_serdes_o0 <= 8'd0;
		main_inout_8x3_serdes_oe <= 1'd0;
		main_inout_8x3_inout_8x3_iinterface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_previous_data <= 1'd0;
		main_inout_8x3_inout_8x3_oe_k <= 1'd0;
		main_inout_8x3_inout_8x3_i_d <= 1'd0;
		main_inout_8x4_serdes_o0 <= 8'd0;
		main_inout_8x4_serdes_oe <= 1'd0;
		main_inout_8x4_inout_8x4_iinterface4_stb <= 1'd0;
		main_inout_8x4_inout_8x4_previous_data <= 1'd0;
		main_inout_8x4_inout_8x4_oe_k <= 1'd0;
		main_inout_8x4_inout_8x4_i_d <= 1'd0;
		main_inout_8x5_serdes_o0 <= 8'd0;
		main_inout_8x5_serdes_oe <= 1'd0;
		main_inout_8x5_inout_8x5_iinterface5_stb <= 1'd0;
		main_inout_8x5_inout_8x5_previous_data <= 1'd0;
		main_inout_8x5_inout_8x5_oe_k <= 1'd0;
		main_inout_8x5_inout_8x5_i_d <= 1'd0;
		main_inout_8x6_serdes_o0 <= 8'd0;
		main_inout_8x6_serdes_oe <= 1'd0;
		main_inout_8x6_inout_8x6_iinterface6_stb <= 1'd0;
		main_inout_8x6_inout_8x6_previous_data <= 1'd0;
		main_inout_8x6_inout_8x6_oe_k <= 1'd0;
		main_inout_8x6_inout_8x6_i_d <= 1'd0;
		main_inout_8x7_serdes_o0 <= 8'd0;
		main_inout_8x7_serdes_oe <= 1'd0;
		main_inout_8x7_inout_8x7_iinterface7_stb <= 1'd0;
		main_inout_8x7_inout_8x7_previous_data <= 1'd0;
		main_inout_8x7_inout_8x7_oe_k <= 1'd0;
		main_inout_8x7_inout_8x7_i_d <= 1'd0;
		main_output_8x0_o <= 8'd0;
		main_output_8x0_previous_data <= 1'd0;
		main_output_8x1_o <= 8'd0;
		main_output_8x1_previous_data <= 1'd0;
		main_output_8x2_o <= 8'd0;
		main_output_8x2_previous_data <= 1'd0;
		main_output_8x3_o <= 8'd0;
		main_output_8x3_previous_data <= 1'd0;
		main_output_8x4_o <= 8'd0;
		main_output_8x4_previous_data <= 1'd0;
		main_output_8x5_o <= 8'd0;
		main_output_8x5_previous_data <= 1'd0;
		main_output_8x6_o <= 8'd0;
		main_output_8x6_previous_data <= 1'd0;
		main_output_8x7_o <= 8'd0;
		main_output_8x7_previous_data <= 1'd0;
		main_spimaster0_interface_cs1 <= 3'd7;
		main_spimaster0_interface_clk <= 1'd0;
		main_spimaster0_spimachine0_cnt <= 7'd0;
		main_spimaster0_spimachine0_do_extend <= 1'd0;
		main_spimaster0_config_offline <= 1'd1;
		main_spimaster0_config_end <= 1'd1;
		main_spimaster0_config_input <= 1'd0;
		main_spimaster0_config_cs_polarity <= 1'd0;
		main_spimaster0_config_clk_polarity <= 1'd0;
		main_spimaster0_config_clk_phase <= 1'd0;
		main_spimaster0_config_lsb_first <= 1'd0;
		main_spimaster0_config_half_duplex <= 1'd0;
		main_spimaster0_config_length <= 5'd0;
		main_spimaster0_config_padding <= 3'd0;
		main_spimaster0_config_div <= 8'd0;
		main_spimaster0_config_cs <= 8'd0;
		main_spimaster0_read <= 1'd0;
		main_output_8x8_o <= 8'd0;
		main_output_8x8_previous_data <= 1'd0;
		main_output_8x9_o <= 8'd0;
		main_output_8x9_previous_data <= 1'd0;
		main_output_8x10_o <= 8'd0;
		main_output_8x10_previous_data <= 1'd0;
		main_output_8x11_o <= 8'd0;
		main_output_8x11_previous_data <= 1'd0;
		main_output_8x12_o <= 8'd0;
		main_output_8x12_previous_data <= 1'd0;
		main_spimaster1_interface_cs1 <= 3'd7;
		main_spimaster1_interface_clk <= 1'd0;
		main_spimaster1_spimachine1_cnt <= 7'd0;
		main_spimaster1_spimachine1_do_extend <= 1'd0;
		main_spimaster1_config_offline <= 1'd1;
		main_spimaster1_config_end <= 1'd1;
		main_spimaster1_config_input <= 1'd0;
		main_spimaster1_config_cs_polarity <= 1'd0;
		main_spimaster1_config_clk_polarity <= 1'd0;
		main_spimaster1_config_clk_phase <= 1'd0;
		main_spimaster1_config_lsb_first <= 1'd0;
		main_spimaster1_config_half_duplex <= 1'd0;
		main_spimaster1_config_length <= 5'd0;
		main_spimaster1_config_padding <= 3'd0;
		main_spimaster1_config_div <= 8'd0;
		main_spimaster1_config_cs <= 8'd0;
		main_spimaster1_read <= 1'd0;
		main_output_8x13_o <= 8'd0;
		main_output_8x13_previous_data <= 1'd0;
		main_output_8x14_o <= 8'd0;
		main_output_8x14_previous_data <= 1'd0;
		main_output_8x15_o <= 8'd0;
		main_output_8x15_previous_data <= 1'd0;
		main_output_8x16_o <= 8'd0;
		main_output_8x16_previous_data <= 1'd0;
		main_output_8x17_o <= 8'd0;
		main_output_8x17_previous_data <= 1'd0;
		main_spimaster2_interface_cs1 <= 3'd7;
		main_spimaster2_interface_clk <= 1'd0;
		main_spimaster2_spimachine2_cnt <= 7'd0;
		main_spimaster2_spimachine2_do_extend <= 1'd0;
		main_spimaster2_config_offline <= 1'd1;
		main_spimaster2_config_end <= 1'd1;
		main_spimaster2_config_input <= 1'd0;
		main_spimaster2_config_cs_polarity <= 1'd0;
		main_spimaster2_config_clk_polarity <= 1'd0;
		main_spimaster2_config_clk_phase <= 1'd0;
		main_spimaster2_config_lsb_first <= 1'd0;
		main_spimaster2_config_half_duplex <= 1'd0;
		main_spimaster2_config_length <= 5'd0;
		main_spimaster2_config_padding <= 3'd0;
		main_spimaster2_config_div <= 8'd0;
		main_spimaster2_config_cs <= 8'd0;
		main_spimaster2_read <= 1'd0;
		main_output_8x18_o <= 8'd0;
		main_output_8x18_previous_data <= 1'd0;
		main_output_8x19_o <= 8'd0;
		main_output_8x19_previous_data <= 1'd0;
		main_output_8x20_o <= 8'd0;
		main_output_8x20_previous_data <= 1'd0;
		main_output_8x21_o <= 8'd0;
		main_output_8x21_previous_data <= 1'd0;
		main_output_8x22_o <= 8'd0;
		main_output_8x22_previous_data <= 1'd0;
		main_output0_pad_k <= 1'd0;
		main_output1_pad_k <= 1'd0;
		builder_spimaster0_state <= 3'd0;
		builder_spimaster1_state <= 3'd0;
		builder_spimaster2_state <= 3'd0;
	end
end

always @(posedge rsys_clk) begin
	main_rtio_core_outputs_lanedistributor_min_minus_timestamp <= (main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp <= (builder_sync_rhs_array_muxed3 - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp <= (builder_sync_rhs_array_muxed4 - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_last_minus_timestamp <= (main_rtio_core_outputs_lanedistributor_last_coarse_timestamp - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_quash <= 1'd0;
	if ((main_rtio_core_cri_chan_sel[15:0] == 6'd36)) begin
		main_rtio_core_outputs_lanedistributor_quash <= 1'd1;
	end
	if (main_rtio_core_outputs_lanedistributor_do_write) begin
		main_rtio_core_outputs_lanedistributor_current_lane <= main_rtio_core_outputs_lanedistributor_use_lanen;
		main_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		builder_sync_t_lhs_array_muxed = main_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		case (main_rtio_core_outputs_lanedistributor_use_lanen)
			1'd0: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= builder_sync_t_lhs_array_muxed;
			end
			1'd1: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= builder_sync_t_lhs_array_muxed;
			end
			2'd2: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= builder_sync_t_lhs_array_muxed;
			end
			2'd3: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= builder_sync_t_lhs_array_muxed;
			end
			3'd4: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= builder_sync_t_lhs_array_muxed;
			end
			3'd5: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= builder_sync_t_lhs_array_muxed;
			end
			3'd6: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= builder_sync_t_lhs_array_muxed;
			end
			default: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= builder_sync_t_lhs_array_muxed;
			end
		endcase
		main_rtio_core_outputs_lanedistributor_seqn <= (main_rtio_core_outputs_lanedistributor_seqn + 1'd1);
	end
	if ((main_rtio_core_cri_cmd == 1'd1)) begin
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
	end
	if (main_rtio_core_outputs_lanedistributor_do_underflow) begin
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd1;
	end
	main_rtio_core_outputs_lanedistributor_sequence_error <= main_rtio_core_outputs_lanedistributor_do_sequence_error;
	main_rtio_core_outputs_lanedistributor_sequence_error_channel <= main_rtio_core_cri_chan_sel[15:0];
	main_rtio_core_outputs_lanedistributor_current_lane_writable_r <= main_rtio_core_outputs_lanedistributor_current_lane_writable;
	if (((~main_rtio_core_outputs_lanedistributor_current_lane_writable_r) & main_rtio_core_outputs_lanedistributor_current_lane_writable)) begin
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd1;
	end
	if (main_rtio_core_outputs_lanedistributor_do_write) begin
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
	end
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
	if ((main_rtio_core_inputs_selected0 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow0 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer0_o) begin
		main_rtio_core_inputs_overflow0 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected1 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow1 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer1_o) begin
		main_rtio_core_inputs_overflow1 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected2 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow2 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer2_o) begin
		main_rtio_core_inputs_overflow2 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected3 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow3 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer3_o) begin
		main_rtio_core_inputs_overflow3 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected4 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow4 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer4_o) begin
		main_rtio_core_inputs_overflow4 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected5 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow5 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer5_o) begin
		main_rtio_core_inputs_overflow5 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected6 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow6 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer6_o) begin
		main_rtio_core_inputs_overflow6 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected7 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow7 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer7_o) begin
		main_rtio_core_inputs_overflow7 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected8 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow8 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer8_o) begin
		main_rtio_core_inputs_overflow8 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected9 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow9 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer9_o) begin
		main_rtio_core_inputs_overflow9 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected10 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow10 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer10_o) begin
		main_rtio_core_inputs_overflow10 <= 1'd1;
	end
	main_rtio_core_inputs_i_ack <= 1'd0;
	if (main_rtio_core_inputs_i_ack) begin
		main_rtio_core_cri_i_status <= {1'd0, main_rtio_core_inputs_i_status_raw[1], (~main_rtio_core_inputs_i_status_raw[0])};
		main_rtio_core_cri_i_data <= builder_sync_t_rhs_array_muxed1;
		main_rtio_core_cri_i_timestamp <= builder_sync_t_rhs_array_muxed2;
	end
	if (((main_rtio_tsc_full_ts_sys >= main_rtio_core_inputs_input_timeout) | (main_rtio_core_inputs_i_status_raw != 1'd0))) begin
		if (main_rtio_core_inputs_input_pending) begin
			main_rtio_core_inputs_i_ack <= 1'd1;
		end
		main_rtio_core_inputs_input_pending <= 1'd0;
	end
	if ((main_rtio_core_cri_cmd == 2'd2)) begin
		main_rtio_core_inputs_input_timeout <= main_rtio_core_cri_i_timeout;
		main_rtio_core_inputs_input_pending <= 1'd1;
		main_rtio_core_cri_i_status <= 3'd4;
	end
	main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
	main_rtio_core_inputs_asyncfifo0_graycounter1_q <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
	main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer0_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer0_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
	main_rtio_core_inputs_asyncfifo1_graycounter3_q <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
	main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer1_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer1_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
	main_rtio_core_inputs_asyncfifo2_graycounter5_q <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
	main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer2_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer2_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
	main_rtio_core_inputs_asyncfifo3_graycounter7_q <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
	main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer3_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer3_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
	main_rtio_core_inputs_asyncfifo4_graycounter9_q <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
	main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer4_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer4_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
	main_rtio_core_inputs_asyncfifo5_graycounter11_q <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
	main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer5_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer5_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
	main_rtio_core_inputs_asyncfifo6_graycounter13_q <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
	main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer6_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer6_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary;
	main_rtio_core_inputs_asyncfifo7_graycounter15_q <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_next;
	main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer7_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer7_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary;
	main_rtio_core_inputs_asyncfifo8_graycounter17_q <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_next;
	main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer8_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer8_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary;
	main_rtio_core_inputs_asyncfifo9_graycounter19_q <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_next;
	main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer9_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer9_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary;
	main_rtio_core_inputs_asyncfifo10_graycounter21_q <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_next;
	main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer10_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer10_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i);
	end
	main_rtio_core_o_collision_sync_ps_toggle_o_r <= main_rtio_core_o_collision_sync_ps_toggle_o;
	if (main_rtio_core_o_collision_sync_ps_ack_i) begin
		main_rtio_core_o_collision_sync_ps_ack_toggle_i <= (~main_rtio_core_o_collision_sync_ps_ack_toggle_i);
	end
	main_rtio_core_o_busy_sync_ps_toggle_o_r <= main_rtio_core_o_busy_sync_ps_toggle_o;
	if (main_rtio_core_o_busy_sync_ps_ack_i) begin
		main_rtio_core_o_busy_sync_ps_ack_toggle_i <= (~main_rtio_core_o_busy_sync_ps_ack_toggle_i);
	end
	if (rsys_rst) begin
		main_rtio_core_cri_i_status <= 4'd0;
		main_rtio_core_outputs_lanedistributor_sequence_error <= 1'd0;
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
		main_rtio_core_outputs_lanedistributor_current_lane <= 3'd0;
		main_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_seqn <= 12'd0;
		main_rtio_core_outputs_lanedistributor_quash <= 1'd0;
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
		main_rtio_core_outputs_lanedistributor_current_lane_writable_r <= 1'd1;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= 8'd0;
		main_rtio_core_inputs_i_ack <= 1'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter1_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow0 <= 1'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter3_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow1 <= 1'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter5_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow2 <= 1'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter7_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow3 <= 1'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter9_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow4 <= 1'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter11_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow5 <= 1'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter13_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow6 <= 1'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter15_q <= 7'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary <= 7'd0;
		main_rtio_core_inputs_overflow7 <= 1'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter17_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary <= 3'd0;
		main_rtio_core_inputs_overflow8 <= 1'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter19_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary <= 3'd0;
		main_rtio_core_inputs_overflow9 <= 1'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter21_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary <= 3'd0;
		main_rtio_core_inputs_overflow10 <= 1'd0;
		main_rtio_core_inputs_input_pending <= 1'd0;
	end
	builder_xilinxmultiregimpl18_regs0 <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q;
	builder_xilinxmultiregimpl18_regs1 <= builder_xilinxmultiregimpl18_regs0;
	builder_xilinxmultiregimpl20_regs0 <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q;
	builder_xilinxmultiregimpl20_regs1 <= builder_xilinxmultiregimpl20_regs0;
	builder_xilinxmultiregimpl22_regs0 <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q;
	builder_xilinxmultiregimpl22_regs1 <= builder_xilinxmultiregimpl22_regs0;
	builder_xilinxmultiregimpl24_regs0 <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q;
	builder_xilinxmultiregimpl24_regs1 <= builder_xilinxmultiregimpl24_regs0;
	builder_xilinxmultiregimpl26_regs0 <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q;
	builder_xilinxmultiregimpl26_regs1 <= builder_xilinxmultiregimpl26_regs0;
	builder_xilinxmultiregimpl28_regs0 <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q;
	builder_xilinxmultiregimpl28_regs1 <= builder_xilinxmultiregimpl28_regs0;
	builder_xilinxmultiregimpl30_regs0 <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q;
	builder_xilinxmultiregimpl30_regs1 <= builder_xilinxmultiregimpl30_regs0;
	builder_xilinxmultiregimpl32_regs0 <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q;
	builder_xilinxmultiregimpl32_regs1 <= builder_xilinxmultiregimpl32_regs0;
	builder_xilinxmultiregimpl33_regs0 <= main_rtio_core_inputs_asyncfifo0_graycounter0_q;
	builder_xilinxmultiregimpl33_regs1 <= builder_xilinxmultiregimpl33_regs0;
	builder_xilinxmultiregimpl35_regs0 <= main_rtio_core_inputs_blindtransfer0_ps_toggle_i;
	builder_xilinxmultiregimpl35_regs1 <= builder_xilinxmultiregimpl35_regs0;
	builder_xilinxmultiregimpl37_regs0 <= main_rtio_core_inputs_asyncfifo1_graycounter2_q;
	builder_xilinxmultiregimpl37_regs1 <= builder_xilinxmultiregimpl37_regs0;
	builder_xilinxmultiregimpl39_regs0 <= main_rtio_core_inputs_blindtransfer1_ps_toggle_i;
	builder_xilinxmultiregimpl39_regs1 <= builder_xilinxmultiregimpl39_regs0;
	builder_xilinxmultiregimpl41_regs0 <= main_rtio_core_inputs_asyncfifo2_graycounter4_q;
	builder_xilinxmultiregimpl41_regs1 <= builder_xilinxmultiregimpl41_regs0;
	builder_xilinxmultiregimpl43_regs0 <= main_rtio_core_inputs_blindtransfer2_ps_toggle_i;
	builder_xilinxmultiregimpl43_regs1 <= builder_xilinxmultiregimpl43_regs0;
	builder_xilinxmultiregimpl45_regs0 <= main_rtio_core_inputs_asyncfifo3_graycounter6_q;
	builder_xilinxmultiregimpl45_regs1 <= builder_xilinxmultiregimpl45_regs0;
	builder_xilinxmultiregimpl47_regs0 <= main_rtio_core_inputs_blindtransfer3_ps_toggle_i;
	builder_xilinxmultiregimpl47_regs1 <= builder_xilinxmultiregimpl47_regs0;
	builder_xilinxmultiregimpl49_regs0 <= main_rtio_core_inputs_asyncfifo4_graycounter8_q;
	builder_xilinxmultiregimpl49_regs1 <= builder_xilinxmultiregimpl49_regs0;
	builder_xilinxmultiregimpl51_regs0 <= main_rtio_core_inputs_blindtransfer4_ps_toggle_i;
	builder_xilinxmultiregimpl51_regs1 <= builder_xilinxmultiregimpl51_regs0;
	builder_xilinxmultiregimpl53_regs0 <= main_rtio_core_inputs_asyncfifo5_graycounter10_q;
	builder_xilinxmultiregimpl53_regs1 <= builder_xilinxmultiregimpl53_regs0;
	builder_xilinxmultiregimpl55_regs0 <= main_rtio_core_inputs_blindtransfer5_ps_toggle_i;
	builder_xilinxmultiregimpl55_regs1 <= builder_xilinxmultiregimpl55_regs0;
	builder_xilinxmultiregimpl57_regs0 <= main_rtio_core_inputs_asyncfifo6_graycounter12_q;
	builder_xilinxmultiregimpl57_regs1 <= builder_xilinxmultiregimpl57_regs0;
	builder_xilinxmultiregimpl59_regs0 <= main_rtio_core_inputs_blindtransfer6_ps_toggle_i;
	builder_xilinxmultiregimpl59_regs1 <= builder_xilinxmultiregimpl59_regs0;
	builder_xilinxmultiregimpl61_regs0 <= main_rtio_core_inputs_asyncfifo7_graycounter14_q;
	builder_xilinxmultiregimpl61_regs1 <= builder_xilinxmultiregimpl61_regs0;
	builder_xilinxmultiregimpl63_regs0 <= main_rtio_core_inputs_blindtransfer7_ps_toggle_i;
	builder_xilinxmultiregimpl63_regs1 <= builder_xilinxmultiregimpl63_regs0;
	builder_xilinxmultiregimpl65_regs0 <= main_rtio_core_inputs_asyncfifo8_graycounter16_q;
	builder_xilinxmultiregimpl65_regs1 <= builder_xilinxmultiregimpl65_regs0;
	builder_xilinxmultiregimpl67_regs0 <= main_rtio_core_inputs_blindtransfer8_ps_toggle_i;
	builder_xilinxmultiregimpl67_regs1 <= builder_xilinxmultiregimpl67_regs0;
	builder_xilinxmultiregimpl69_regs0 <= main_rtio_core_inputs_asyncfifo9_graycounter18_q;
	builder_xilinxmultiregimpl69_regs1 <= builder_xilinxmultiregimpl69_regs0;
	builder_xilinxmultiregimpl71_regs0 <= main_rtio_core_inputs_blindtransfer9_ps_toggle_i;
	builder_xilinxmultiregimpl71_regs1 <= builder_xilinxmultiregimpl71_regs0;
	builder_xilinxmultiregimpl73_regs0 <= main_rtio_core_inputs_asyncfifo10_graycounter20_q;
	builder_xilinxmultiregimpl73_regs1 <= builder_xilinxmultiregimpl73_regs0;
	builder_xilinxmultiregimpl75_regs0 <= main_rtio_core_inputs_blindtransfer10_ps_toggle_i;
	builder_xilinxmultiregimpl75_regs1 <= builder_xilinxmultiregimpl75_regs0;
	builder_xilinxmultiregimpl77_regs0 <= main_rtio_core_o_collision_sync_ps_toggle_i;
	builder_xilinxmultiregimpl77_regs1 <= builder_xilinxmultiregimpl77_regs0;
	builder_xilinxmultiregimpl79_regs0 <= main_rtio_core_o_collision_sync_bxfer_data;
	builder_xilinxmultiregimpl79_regs1 <= builder_xilinxmultiregimpl79_regs0;
	builder_xilinxmultiregimpl80_regs0 <= main_rtio_core_o_busy_sync_ps_toggle_i;
	builder_xilinxmultiregimpl80_regs1 <= builder_xilinxmultiregimpl80_regs0;
	builder_xilinxmultiregimpl82_regs0 <= main_rtio_core_o_busy_sync_bxfer_data;
	builder_xilinxmultiregimpl82_regs1 <= builder_xilinxmultiregimpl82_regs0;
end

always @(posedge rtio_clk) begin
	if (main_rtio_tsc_load) begin
		main_rtio_tsc_coarse_ts <= main_rtio_tsc_load_value;
	end else begin
		main_rtio_tsc_coarse_ts <= (main_rtio_tsc_coarse_ts + 1'd1);
	end
	main_rtio_tsc_value_gray_rtio <= (main_rtio_tsc_i ^ main_rtio_tsc_i[60:1]);
	if (rtio_rst) begin
		main_rtio_tsc_coarse_ts <= 61'd0;
	end
end

always @(posedge sys_clk) begin
	main_genericstandalone_genericstandalone_genericstandalone_tmpu_error <= 1'd0;
	if ((main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage & (main_genericstandalone_genericstandalone_genericstandalone_dbus_adr[29:10] == 1'd0))) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_error <= 1'd1;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage & (main_genericstandalone_genericstandalone_genericstandalone_dbus_adr[29:10] == main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage))) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_error <= 1'd1;
	end
	main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd0;
	if (((main_genericstandalone_genericstandalone_genericstandalone_sram_bus_cyc & main_genericstandalone_genericstandalone_genericstandalone_sram_bus_stb) & (~main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack))) begin
		main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd1;
	end
	main_genericstandalone_genericstandalone_genericstandalone_interface_we <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_w;
	main_genericstandalone_genericstandalone_genericstandalone_interface_adr <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_adr;
	main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_interface_dat_r;
	if ((main_genericstandalone_genericstandalone_genericstandalone_counter == 1'd1)) begin
		main_genericstandalone_genericstandalone_genericstandalone_interface_we <= main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_we;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_counter == 2'd2)) begin
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd1;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_counter == 2'd3)) begin
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_genericstandalone_counter != 1'd0)) begin
		main_genericstandalone_genericstandalone_genericstandalone_counter <= (main_genericstandalone_genericstandalone_genericstandalone_counter + 1'd1);
	end else begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_cyc & main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_stb)) begin
			main_genericstandalone_genericstandalone_genericstandalone_counter <= 1'd1;
		end
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd0;
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_stb & (~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy)) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_payload_data;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen & main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount + 1'd1);
			if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd0;
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd1;
				end else begin
					serial_tx <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg[0];
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= {1'd0, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy) begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx} <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx + main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage);
	end else begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd0;
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx;
	if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy)) begin
		if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) & main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd1;
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount + 1'd1);
			if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount == 1'd0)) begin
				if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount == 4'd9)) begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
					if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx) begin
						main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data <= main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg;
						main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd1;
					end
				end else begin
					main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg <= {main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy) begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx} <= (main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx + main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage);
	end else begin
		{main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen, main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_trigger) & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd1;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_trigger) & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd1;
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_replace))) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_do_read) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace))) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_we & main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_syncfifo_writable) & (~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_replace))) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read)) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_do_read) begin
			main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level - 1'd1);
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage) begin
		if ((main_genericstandalone_genericstandalone_genericstandalone_timer0_value == 1'd0)) begin
			main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage;
		end else begin
			main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= (main_genericstandalone_genericstandalone_genericstandalone_timer0_value - 1'd1);
		end
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status <= main_genericstandalone_genericstandalone_genericstandalone_timer0_value;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_clear) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd0;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger <= main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger;
	if (((~main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_trigger) & main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger)) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd1;
	end
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 <= main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_en;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2;
	main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid <= main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4;
	main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en <= {main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en[2:0], main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_en};
	main_genericstandalone_genericstandalone_ddrphy_oe_dqs <= main_genericstandalone_genericstandalone_ddrphy_oe;
	main_genericstandalone_genericstandalone_ddrphy_oe_dq <= main_genericstandalone_genericstandalone_ddrphy_oe;
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p0_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p1_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p2_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata_valid) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status <= main_genericstandalone_genericstandalone_genericstandalone_inti_p3_rddata;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce0) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset0) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce1) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset1) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce2) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset2) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce3) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset3) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce4) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset4) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce5) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset5) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce6) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset6) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_ce7) begin
		if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_open) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd0;
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row0;
		end
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_reset7) begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= 15'd0;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_wait) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_done)) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count <= (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count - 1'd1);
		end
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count <= 3'd4;
	end
	if (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_wait) begin
		if ((~main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_done)) begin
			main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count <= (main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count - 1'd1);
		end
	end else begin
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count <= 10'd886;
	end
	builder_minicon_state <= builder_minicon_next_state;
	main_genericstandalone_genericstandalone_genericstandalone_adr_offset_r <= main_genericstandalone_genericstandalone_genericstandalone_cpulevel_sdram_if_arbitrated_adr[1:0];
	builder_fullmemorywe_state <= builder_fullmemorywe_next_state;
	if ((main_genericstandalone_genericstandalone_spiflash_i1 == 1'd0)) begin
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_dqi <= main_genericstandalone_genericstandalone_spiflash_i0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1)) begin
		main_genericstandalone_genericstandalone_spiflash_i1 <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr <= {main_genericstandalone_genericstandalone_spiflash_sr[29:0], main_genericstandalone_genericstandalone_spiflash_dqi};
	end else begin
		main_genericstandalone_genericstandalone_spiflash_i1 <= (main_genericstandalone_genericstandalone_spiflash_i1 + 1'd1);
	end
	if ((((main_genericstandalone_genericstandalone_spiflash_bus_cyc & main_genericstandalone_genericstandalone_spiflash_bus_stb) & (main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1)) & (main_genericstandalone_genericstandalone_spiflash_counter == 1'd0))) begin
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr[31:16] <= 16'd61423;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 5'd16)) begin
		main_genericstandalone_genericstandalone_spiflash_sr[31:8] <= {main_genericstandalone_genericstandalone_spiflash_bus_adr, {2{1'd0}}};
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 6'd40)) begin
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 7'd82)) begin
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd1;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 7'd83)) begin
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd0;
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 7'd85)) begin
	end
	if ((main_genericstandalone_genericstandalone_spiflash_counter == 7'd85)) begin
		main_genericstandalone_genericstandalone_spiflash_counter <= 1'd0;
	end else begin
		if ((main_genericstandalone_genericstandalone_spiflash_counter != 1'd0)) begin
			main_genericstandalone_genericstandalone_spiflash_counter <= (main_genericstandalone_genericstandalone_spiflash_counter + 1'd1);
		end else begin
			if (((main_genericstandalone_genericstandalone_spiflash_bus_cyc & main_genericstandalone_genericstandalone_spiflash_bus_stb) & (main_genericstandalone_genericstandalone_spiflash_i1 == 1'd1))) begin
				main_genericstandalone_genericstandalone_spiflash_counter <= 1'd1;
			end
		end
	end
	main_genericstandalone_tx_mmcm_reset <= (~main_genericstandalone_genericstandalone_qpll_lock);
	if (main_genericstandalone_rx_reset) begin
		main_genericstandalone_cdr_locked <= 1'd0;
		main_genericstandalone_cdr_lock_counter <= 1'd0;
	end else begin
		if ((main_genericstandalone_cdr_lock_counter != 13'd4531)) begin
			main_genericstandalone_cdr_lock_counter <= (main_genericstandalone_cdr_lock_counter + 1'd1);
		end else begin
			main_genericstandalone_cdr_locked <= 1'd1;
		end
	end
	main_genericstandalone_rx_mmcm_reset <= (~main_genericstandalone_cdr_locked);
	main_genericstandalone_tx_init_qpll_reset0 <= main_genericstandalone_tx_init_qpll_reset1;
	main_genericstandalone_tx_init_tx_reset0 <= main_genericstandalone_tx_init_tx_reset1;
	main_genericstandalone_tx_init_tick <= 1'd0;
	if ((main_genericstandalone_tx_init_timer == 6'd57)) begin
		main_genericstandalone_tx_init_tick <= 1'd1;
		main_genericstandalone_tx_init_timer <= 1'd0;
	end else begin
		main_genericstandalone_tx_init_timer <= (main_genericstandalone_tx_init_timer + 1'd1);
	end
	builder_a7_1000basex_gtptxinit_state <= builder_a7_1000basex_gtptxinit_next_state;
	main_genericstandalone_rx_init_rx_reset0 <= main_genericstandalone_rx_init_rx_reset1;
	main_genericstandalone_rx_init_rx_pma_reset_done_r <= main_genericstandalone_rx_init_rx_pma_reset_done1;
	builder_a7_1000basex_gtprxinit_state <= builder_a7_1000basex_gtprxinit_next_state;
	if (main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value_ce) begin
		main_genericstandalone_rx_init_drpvalue <= main_genericstandalone_rx_init_drpvalue_gtprxinit_next_value;
	end
	main_genericstandalone_toggle_o_r <= main_genericstandalone_toggle_o;
	if (main_genericstandalone_ps_preamble_error_o) begin
		main_genericstandalone_preamble_errors_status <= (main_genericstandalone_preamble_errors_status + 1'd1);
	end
	if (main_genericstandalone_ps_crc_error_o) begin
		main_genericstandalone_crc_errors_status <= (main_genericstandalone_crc_errors_status + 1'd1);
	end
	main_genericstandalone_ps_preamble_error_toggle_o_r <= main_genericstandalone_ps_preamble_error_toggle_o;
	main_genericstandalone_ps_crc_error_toggle_o_r <= main_genericstandalone_ps_crc_error_toggle_o;
	main_genericstandalone_tx_cdc_graycounter0_q_binary <= main_genericstandalone_tx_cdc_graycounter0_q_next_binary;
	main_genericstandalone_tx_cdc_graycounter0_q <= main_genericstandalone_tx_cdc_graycounter0_q_next;
	main_genericstandalone_rx_cdc_graycounter1_q_binary <= main_genericstandalone_rx_cdc_graycounter1_q_next_binary;
	main_genericstandalone_rx_cdc_graycounter1_q <= main_genericstandalone_rx_cdc_graycounter1_q_next;
	if (main_genericstandalone_writer_counter_reset) begin
		main_genericstandalone_writer_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_writer_counter_ce) begin
			main_genericstandalone_writer_counter <= (main_genericstandalone_writer_counter + main_genericstandalone_writer_increment);
		end
	end
	if (main_genericstandalone_writer_slot_ce) begin
		main_genericstandalone_writer_slot <= (main_genericstandalone_writer_slot + 1'd1);
	end
	if (((main_genericstandalone_writer_fifo_syncfifo_we & main_genericstandalone_writer_fifo_syncfifo_writable) & (~main_genericstandalone_writer_fifo_replace))) begin
		main_genericstandalone_writer_fifo_produce <= (main_genericstandalone_writer_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_writer_fifo_do_read) begin
		main_genericstandalone_writer_fifo_consume <= (main_genericstandalone_writer_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_writer_fifo_syncfifo_we & main_genericstandalone_writer_fifo_syncfifo_writable) & (~main_genericstandalone_writer_fifo_replace))) begin
		if ((~main_genericstandalone_writer_fifo_do_read)) begin
			main_genericstandalone_writer_fifo_level <= (main_genericstandalone_writer_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_writer_fifo_do_read) begin
			main_genericstandalone_writer_fifo_level <= (main_genericstandalone_writer_fifo_level - 1'd1);
		end
	end
	builder_liteethmacsramwriter_state <= builder_liteethmacsramwriter_next_state;
	if (main_genericstandalone_writer_errors_status_next_value_ce) begin
		main_genericstandalone_writer_errors_status <= main_genericstandalone_writer_errors_status_next_value;
	end
	if (main_genericstandalone_reader_counter_reset) begin
		main_genericstandalone_reader_counter <= 1'd0;
	end else begin
		if (main_genericstandalone_reader_counter_ce) begin
			main_genericstandalone_reader_counter <= (main_genericstandalone_reader_counter + 3'd4);
		end
	end
	main_genericstandalone_reader_last_d <= main_genericstandalone_reader_last;
	if (main_genericstandalone_reader_done_clear) begin
		main_genericstandalone_reader_done_pending <= 1'd0;
	end
	if (main_genericstandalone_reader_done_trigger) begin
		main_genericstandalone_reader_done_pending <= 1'd1;
	end
	if (((main_genericstandalone_reader_fifo_syncfifo_we & main_genericstandalone_reader_fifo_syncfifo_writable) & (~main_genericstandalone_reader_fifo_replace))) begin
		main_genericstandalone_reader_fifo_produce <= (main_genericstandalone_reader_fifo_produce + 1'd1);
	end
	if (main_genericstandalone_reader_fifo_do_read) begin
		main_genericstandalone_reader_fifo_consume <= (main_genericstandalone_reader_fifo_consume + 1'd1);
	end
	if (((main_genericstandalone_reader_fifo_syncfifo_we & main_genericstandalone_reader_fifo_syncfifo_writable) & (~main_genericstandalone_reader_fifo_replace))) begin
		if ((~main_genericstandalone_reader_fifo_do_read)) begin
			main_genericstandalone_reader_fifo_level <= (main_genericstandalone_reader_fifo_level + 1'd1);
		end
	end else begin
		if (main_genericstandalone_reader_fifo_do_read) begin
			main_genericstandalone_reader_fifo_level <= (main_genericstandalone_reader_fifo_level - 1'd1);
		end
	end
	builder_liteethmacsramreader_state <= builder_liteethmacsramreader_next_state;
	main_genericstandalone_sram0_bus_ack0 <= 1'd0;
	if (((main_genericstandalone_sram0_bus_cyc0 & main_genericstandalone_sram0_bus_stb0) & (~main_genericstandalone_sram0_bus_ack0))) begin
		main_genericstandalone_sram0_bus_ack0 <= 1'd1;
	end
	main_genericstandalone_sram1_bus_ack0 <= 1'd0;
	if (((main_genericstandalone_sram1_bus_cyc0 & main_genericstandalone_sram1_bus_stb0) & (~main_genericstandalone_sram1_bus_ack0))) begin
		main_genericstandalone_sram1_bus_ack0 <= 1'd1;
	end
	main_genericstandalone_sram2_bus_ack0 <= 1'd0;
	if (((main_genericstandalone_sram2_bus_cyc0 & main_genericstandalone_sram2_bus_stb0) & (~main_genericstandalone_sram2_bus_ack0))) begin
		main_genericstandalone_sram2_bus_ack0 <= 1'd1;
	end
	main_genericstandalone_sram3_bus_ack0 <= 1'd0;
	if (((main_genericstandalone_sram3_bus_cyc0 & main_genericstandalone_sram3_bus_stb0) & (~main_genericstandalone_sram3_bus_ack0))) begin
		main_genericstandalone_sram3_bus_ack0 <= 1'd1;
	end
	main_genericstandalone_sram0_bus_ack1 <= 1'd0;
	if (((main_genericstandalone_sram0_bus_cyc1 & main_genericstandalone_sram0_bus_stb1) & (~main_genericstandalone_sram0_bus_ack1))) begin
		main_genericstandalone_sram0_bus_ack1 <= 1'd1;
	end
	main_genericstandalone_sram1_bus_ack1 <= 1'd0;
	if (((main_genericstandalone_sram1_bus_cyc1 & main_genericstandalone_sram1_bus_stb1) & (~main_genericstandalone_sram1_bus_ack1))) begin
		main_genericstandalone_sram1_bus_ack1 <= 1'd1;
	end
	main_genericstandalone_sram2_bus_ack1 <= 1'd0;
	if (((main_genericstandalone_sram2_bus_cyc1 & main_genericstandalone_sram2_bus_stb1) & (~main_genericstandalone_sram2_bus_ack1))) begin
		main_genericstandalone_sram2_bus_ack1 <= 1'd1;
	end
	main_genericstandalone_sram3_bus_ack1 <= 1'd0;
	if (((main_genericstandalone_sram3_bus_cyc1 & main_genericstandalone_sram3_bus_stb1) & (~main_genericstandalone_sram3_bus_ack1))) begin
		main_genericstandalone_sram3_bus_ack1 <= 1'd1;
	end
	main_genericstandalone_slave_sel_r <= main_genericstandalone_slave_sel;
	case (builder_grant)
		1'd0: begin
			if ((~builder_request[0])) begin
				if (builder_request[1]) begin
					builder_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_request[1])) begin
				if (builder_request[0]) begin
					builder_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_slave_sel_r <= builder_slave_sel;
	main_genericstandalone_mailbox_i1_dat_r <= builder_sync_rhs_array_muxed5;
	main_genericstandalone_mailbox_i1_ack <= 1'd0;
	if (((main_genericstandalone_mailbox_i1_cyc & main_genericstandalone_mailbox_i1_stb) & (~main_genericstandalone_mailbox_i1_ack))) begin
		main_genericstandalone_mailbox_i1_ack <= 1'd1;
		if (main_genericstandalone_mailbox_i1_we) begin
			builder_sync_t_t_array_muxed0 = main_genericstandalone_mailbox_i1_dat_w;
			case (main_genericstandalone_mailbox_i1_adr[1:0])
				1'd0: begin
					main_genericstandalone_mailbox0 <= builder_sync_t_t_array_muxed0;
				end
				1'd1: begin
					main_genericstandalone_mailbox1 <= builder_sync_t_t_array_muxed0;
				end
				default: begin
					main_genericstandalone_mailbox2 <= builder_sync_t_t_array_muxed0;
				end
			endcase
		end
	end
	main_genericstandalone_mailbox_i2_dat_r <= builder_sync_rhs_array_muxed6;
	main_genericstandalone_mailbox_i2_ack <= 1'd0;
	if (((main_genericstandalone_mailbox_i2_cyc & main_genericstandalone_mailbox_i2_stb) & (~main_genericstandalone_mailbox_i2_ack))) begin
		main_genericstandalone_mailbox_i2_ack <= 1'd1;
		if (main_genericstandalone_mailbox_i2_we) begin
			builder_sync_t_t_array_muxed1 = main_genericstandalone_mailbox_i2_dat_w;
			case (main_genericstandalone_mailbox_i2_adr[1:0])
				1'd0: begin
					main_genericstandalone_mailbox0 <= builder_sync_t_t_array_muxed1;
				end
				1'd1: begin
					main_genericstandalone_mailbox1 <= builder_sync_t_t_array_muxed1;
				end
				default: begin
					main_genericstandalone_mailbox2 <= builder_sync_t_t_array_muxed1;
				end
			endcase
		end
	end
	main_rtio_tsc_o <= main_rtio_tsc_value_sys;
	main_rtio_core_cmd_reset <= main_rtio_core_reset_re;
	main_rtio_core_cmd_reset_phy <= main_rtio_core_reset_phy_re;
	main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= (main_rtio_tsc_coarse_ts_sys + 5'd16);
	if (main_rtio_core_async_error_re) begin
		if (main_rtio_core_async_error_r[0]) begin
			main_rtio_core_o_collision <= 1'd0;
		end
		if (main_rtio_core_async_error_r[1]) begin
			main_rtio_core_o_busy <= 1'd0;
		end
		if (main_rtio_core_async_error_r[2]) begin
			main_rtio_core_o_sequence_error <= 1'd0;
		end
	end
	if (main_rtio_core_o_collision_sync_o) begin
		main_rtio_core_o_collision <= 1'd1;
		if ((~main_rtio_core_o_collision)) begin
			main_rtio_core_collision_channel_status <= main_rtio_core_o_collision_sync_data_o;
		end
	end
	if (main_rtio_core_o_busy_sync_o) begin
		main_rtio_core_o_busy <= 1'd1;
		if ((~main_rtio_core_o_busy)) begin
			main_rtio_core_busy_channel_status <= main_rtio_core_o_busy_sync_data_o;
		end
	end
	if (main_rtio_core_outputs_lanedistributor_sequence_error) begin
		main_rtio_core_o_sequence_error <= 1'd1;
		if ((~main_rtio_core_o_sequence_error)) begin
			main_rtio_core_sequence_error_channel_status <= main_rtio_core_outputs_lanedistributor_sequence_error_channel;
		end
	end
	if (main_rtio_now_hi_re) begin
		main_rtio_now_hi_backing <= main_rtio_now_hi_r;
	end
	if (main_rtio_now_lo_re) begin
		main_rtio_now <= {main_rtio_now_hi_backing, main_rtio_now_lo_r};
	end
	if (main_rtio_counter_update_re) begin
		main_rtio_counter_status <= main_rtio_tsc_full_ts_sys;
	end
	case (main_genericstandalone_csrbank0_bus_adr[4:0])
		1'd0: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_target0_w;
		end
		1'd1: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_rtio_now_hi_w;
		end
		2'd2: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_rtio_now_lo_w;
		end
		2'd3: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data15_w;
		end
		3'd4: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data14_w;
		end
		3'd5: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data13_w;
		end
		3'd6: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data12_w;
		end
		3'd7: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data11_w;
		end
		4'd8: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data10_w;
		end
		4'd9: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data9_w;
		end
		4'd10: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data8_w;
		end
		4'd11: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data7_w;
		end
		4'd12: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data6_w;
		end
		4'd13: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data5_w;
		end
		4'd14: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data4_w;
		end
		4'd15: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data3_w;
		end
		5'd16: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data2_w;
		end
		5'd17: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data1_w;
		end
		5'd18: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_data0_w;
		end
		5'd19: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_o_status_w;
		end
		5'd20: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_timeout1_w;
		end
		5'd21: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_timeout0_w;
		end
		5'd22: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_data_w;
		end
		5'd23: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_timestamp1_w;
		end
		5'd24: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_timestamp0_w;
		end
		5'd25: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_i_status_w;
		end
		5'd26: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_rtio_i_overflow_reset_w;
		end
		5'd27: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_counter1_w;
		end
		5'd28: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_genericstandalone_csrbank0_counter0_w;
		end
		5'd29: begin
			main_genericstandalone_csrbank0_bus_dat_r <= main_rtio_counter_update_w;
		end
	endcase
	if (main_genericstandalone_csrbank0_bus_ack) begin
		main_genericstandalone_csrbank0_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_csrbank0_bus_cyc & main_genericstandalone_csrbank0_bus_stb)) begin
			main_genericstandalone_csrbank0_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_csrbank0_target0_re) begin
		main_rtio_target_storage_full[31:0] <= main_genericstandalone_csrbank0_target0_r;
	end
	main_rtio_target_re <= main_genericstandalone_csrbank0_target0_re;
	if (main_rtio_o_data_we) begin
		main_rtio_o_data_storage_full <= (main_rtio_o_data_dat_w <<< 1'd0);
	end
	if (main_genericstandalone_csrbank0_o_data15_re) begin
		main_rtio_o_data_storage_full[511:480] <= main_genericstandalone_csrbank0_o_data15_r;
	end
	if (main_genericstandalone_csrbank0_o_data14_re) begin
		main_rtio_o_data_storage_full[479:448] <= main_genericstandalone_csrbank0_o_data14_r;
	end
	if (main_genericstandalone_csrbank0_o_data13_re) begin
		main_rtio_o_data_storage_full[447:416] <= main_genericstandalone_csrbank0_o_data13_r;
	end
	if (main_genericstandalone_csrbank0_o_data12_re) begin
		main_rtio_o_data_storage_full[415:384] <= main_genericstandalone_csrbank0_o_data12_r;
	end
	if (main_genericstandalone_csrbank0_o_data11_re) begin
		main_rtio_o_data_storage_full[383:352] <= main_genericstandalone_csrbank0_o_data11_r;
	end
	if (main_genericstandalone_csrbank0_o_data10_re) begin
		main_rtio_o_data_storage_full[351:320] <= main_genericstandalone_csrbank0_o_data10_r;
	end
	if (main_genericstandalone_csrbank0_o_data9_re) begin
		main_rtio_o_data_storage_full[319:288] <= main_genericstandalone_csrbank0_o_data9_r;
	end
	if (main_genericstandalone_csrbank0_o_data8_re) begin
		main_rtio_o_data_storage_full[287:256] <= main_genericstandalone_csrbank0_o_data8_r;
	end
	if (main_genericstandalone_csrbank0_o_data7_re) begin
		main_rtio_o_data_storage_full[255:224] <= main_genericstandalone_csrbank0_o_data7_r;
	end
	if (main_genericstandalone_csrbank0_o_data6_re) begin
		main_rtio_o_data_storage_full[223:192] <= main_genericstandalone_csrbank0_o_data6_r;
	end
	if (main_genericstandalone_csrbank0_o_data5_re) begin
		main_rtio_o_data_storage_full[191:160] <= main_genericstandalone_csrbank0_o_data5_r;
	end
	if (main_genericstandalone_csrbank0_o_data4_re) begin
		main_rtio_o_data_storage_full[159:128] <= main_genericstandalone_csrbank0_o_data4_r;
	end
	if (main_genericstandalone_csrbank0_o_data3_re) begin
		main_rtio_o_data_storage_full[127:96] <= main_genericstandalone_csrbank0_o_data3_r;
	end
	if (main_genericstandalone_csrbank0_o_data2_re) begin
		main_rtio_o_data_storage_full[95:64] <= main_genericstandalone_csrbank0_o_data2_r;
	end
	if (main_genericstandalone_csrbank0_o_data1_re) begin
		main_rtio_o_data_storage_full[63:32] <= main_genericstandalone_csrbank0_o_data1_r;
	end
	if (main_genericstandalone_csrbank0_o_data0_re) begin
		main_rtio_o_data_storage_full[31:0] <= main_genericstandalone_csrbank0_o_data0_r;
	end
	main_rtio_o_data_re <= main_genericstandalone_csrbank0_o_data0_re;
	if (main_genericstandalone_csrbank0_i_timeout1_re) begin
		main_rtio_i_timeout_storage_full[63:32] <= main_genericstandalone_csrbank0_i_timeout1_r;
	end
	if (main_genericstandalone_csrbank0_i_timeout0_re) begin
		main_rtio_i_timeout_storage_full[31:0] <= main_genericstandalone_csrbank0_i_timeout0_r;
	end
	main_rtio_i_timeout_re <= main_genericstandalone_csrbank0_i_timeout0_re;
	case (main_genericstandalone_csrbank1_bus_adr[3:0])
		1'd0: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_dma_enable_enable_w;
		end
		1'd1: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_base_address1_w;
		end
		2'd2: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_base_address0_w;
		end
		2'd3: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_time_offset1_w;
		end
		3'd4: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_time_offset0_w;
		end
		3'd5: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_dma_cri_master_error_w;
		end
		3'd6: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_error_channel_w;
		end
		3'd7: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_error_timestamp1_w;
		end
		4'd8: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_error_timestamp0_w;
		end
		4'd9: begin
			main_genericstandalone_csrbank1_bus_dat_r <= main_genericstandalone_csrbank1_error_address_w;
		end
	endcase
	if (main_genericstandalone_csrbank1_bus_ack) begin
		main_genericstandalone_csrbank1_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_csrbank1_bus_cyc & main_genericstandalone_csrbank1_bus_stb)) begin
			main_genericstandalone_csrbank1_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_csrbank1_base_address1_re) begin
		main_dma_dma_storage_full[33:32] <= main_genericstandalone_csrbank1_base_address1_r;
	end
	if (main_genericstandalone_csrbank1_base_address0_re) begin
		main_dma_dma_storage_full[31:0] <= main_genericstandalone_csrbank1_base_address0_r;
	end
	main_dma_dma_re <= main_genericstandalone_csrbank1_base_address0_re;
	if (main_genericstandalone_csrbank1_time_offset1_re) begin
		main_dma_time_offset_storage_full[63:32] <= main_genericstandalone_csrbank1_time_offset1_r;
	end
	if (main_genericstandalone_csrbank1_time_offset0_re) begin
		main_dma_time_offset_storage_full[31:0] <= main_genericstandalone_csrbank1_time_offset0_r;
	end
	main_dma_time_offset_re <= main_genericstandalone_csrbank1_time_offset0_re;
	main_cri_con_selected <= main_cri_con_shared_chan_sel[23:16];
	case (main_genericstandalone_csrbank2_bus_adr[0])
		1'd0: begin
			main_genericstandalone_csrbank2_bus_dat_r <= main_genericstandalone_csrbank2_selected0_w;
		end
	endcase
	if (main_genericstandalone_csrbank2_bus_ack) begin
		main_genericstandalone_csrbank2_bus_ack <= 1'd0;
	end else begin
		if ((main_genericstandalone_csrbank2_bus_cyc & main_genericstandalone_csrbank2_bus_stb)) begin
			main_genericstandalone_csrbank2_bus_ack <= 1'd1;
		end
	end
	if (main_genericstandalone_csrbank2_selected0_re) begin
		main_cri_con_storage_full[1:0] <= main_genericstandalone_csrbank2_selected0_r;
	end
	main_cri_con_re <= main_genericstandalone_csrbank2_selected0_re;
	if (main_mon_value_update_re) begin
		main_mon_status <= builder_sync_t_rhs_array_muxed3;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd0)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys0 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd0)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys1 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd0)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys2 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd1)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys3 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd1)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys4 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd1)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys5 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd2)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys6 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd2)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys7 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd2)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys8 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys9 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys10 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys11 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd4)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys12 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd4)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys13 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd4)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys14 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd5)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys15 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd5)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys16 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd5)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys17 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd6)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys18 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd6)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys19 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd6)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys20 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys21 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys22 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys23 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd8)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys24 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd8)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys25 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd9)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys26 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd9)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys27 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd10)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys28 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd10)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys29 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd11)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys30 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd11)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys31 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd12)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys32 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd12)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys33 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd13)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys34 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd13)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys35 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd14)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys36 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd14)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys37 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd15)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys38 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd15)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys39 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd17)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys40 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd17)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys41 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd18)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys42 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd18)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys43 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd19)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys44 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd19)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys45 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd20)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys46 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd20)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys47 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd21)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys48 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd21)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys49 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd23)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys50 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd23)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys51 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd24)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys52 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd24)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys53 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd25)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys54 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd25)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys55 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd26)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys56 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd26)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys57 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd27)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys58 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd27)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys59 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd29)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys60 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd29)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys61 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd30)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys62 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd30)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys63 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd31)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys64 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd31)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys65 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd32)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys66 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd32)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys67 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd33)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys68 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd33)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys69 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd34)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys70 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd34)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys71 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd35)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys72 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 6'd35)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys73 <= main_inj_value_r;
	end
	main_rtio_analyzer_enable_r <= main_rtio_analyzer_enable_storage;
	if ((main_rtio_analyzer_enable_storage & (~main_rtio_analyzer_enable_r))) begin
		main_rtio_analyzer_busy_status <= 1'd1;
	end
	if (((main_rtio_analyzer_dma_sink_stb & main_rtio_analyzer_dma_sink_ack) & main_rtio_analyzer_dma_sink_eop)) begin
		main_rtio_analyzer_busy_status <= 1'd0;
	end
	main_rtio_analyzer_message_encoder_read_wait_event_r <= main_rtio_core_cri_i_status[2];
	main_rtio_analyzer_message_encoder_just_written <= (main_rtio_core_cri_cmd == 1'd1);
	main_rtio_analyzer_message_encoder_enable_r <= main_rtio_analyzer_enable_storage;
	if (((~main_rtio_analyzer_enable_storage) & main_rtio_analyzer_message_encoder_enable_r)) begin
		main_rtio_analyzer_message_encoder_stopping <= 1'd1;
	end
	if ((~main_rtio_analyzer_message_encoder_stopping)) begin
		if (main_rtio_analyzer_message_encoder_exception_stb) begin
			main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_exception_padding1, main_rtio_analyzer_message_encoder_exception_exception_type, main_rtio_analyzer_message_encoder_exception_rtio_counter, main_rtio_analyzer_message_encoder_exception_padding0, main_rtio_analyzer_message_encoder_exception_channel, main_rtio_analyzer_message_encoder_exception_message_type};
		end else begin
			main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_input_output_data, main_rtio_analyzer_message_encoder_input_output_address_padding, main_rtio_analyzer_message_encoder_input_output_rtio_counter, main_rtio_analyzer_message_encoder_input_output_timestamp, main_rtio_analyzer_message_encoder_input_output_channel, main_rtio_analyzer_message_encoder_input_output_message_type};
		end
		main_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_rtio_analyzer_message_encoder_source_stb <= (main_rtio_analyzer_enable_storage & (main_rtio_analyzer_message_encoder_input_output_stb | main_rtio_analyzer_message_encoder_exception_stb));
		if (main_rtio_analyzer_message_encoder_overflow_reset_re) begin
			main_rtio_analyzer_message_encoder_status <= 1'd0;
		end
		if ((main_rtio_analyzer_message_encoder_source_stb & (~main_rtio_analyzer_message_encoder_source_ack))) begin
			main_rtio_analyzer_message_encoder_status <= 1'd1;
		end
	end else begin
		main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_stopped_padding1, main_rtio_analyzer_message_encoder_stopped_rtio_counter, main_rtio_analyzer_message_encoder_stopped_padding0, main_rtio_analyzer_message_encoder_stopped_message_type};
		main_rtio_analyzer_message_encoder_source_eop <= 1'd1;
		main_rtio_analyzer_message_encoder_source_stb <= 1'd1;
		if (main_rtio_analyzer_message_encoder_source_ack) begin
			main_rtio_analyzer_message_encoder_stopping <= 1'd0;
		end
	end
	if (main_rtio_analyzer_fifo_syncfifo_re) begin
		main_rtio_analyzer_fifo_readable <= 1'd1;
	end else begin
		if (main_rtio_analyzer_fifo_re) begin
			main_rtio_analyzer_fifo_readable <= 1'd0;
		end
	end
	if (((main_rtio_analyzer_fifo_syncfifo_we & main_rtio_analyzer_fifo_syncfifo_writable) & (~main_rtio_analyzer_fifo_replace))) begin
		main_rtio_analyzer_fifo_produce <= (main_rtio_analyzer_fifo_produce + 1'd1);
	end
	if (main_rtio_analyzer_fifo_do_read) begin
		main_rtio_analyzer_fifo_consume <= (main_rtio_analyzer_fifo_consume + 1'd1);
	end
	if (((main_rtio_analyzer_fifo_syncfifo_we & main_rtio_analyzer_fifo_syncfifo_writable) & (~main_rtio_analyzer_fifo_replace))) begin
		if ((~main_rtio_analyzer_fifo_do_read)) begin
			main_rtio_analyzer_fifo_level0 <= (main_rtio_analyzer_fifo_level0 + 1'd1);
		end
	end else begin
		if (main_rtio_analyzer_fifo_do_read) begin
			main_rtio_analyzer_fifo_level0 <= (main_rtio_analyzer_fifo_level0 - 1'd1);
		end
	end
	if ((main_rtio_analyzer_converter_source_stb & main_rtio_analyzer_converter_source_ack)) begin
		if (main_rtio_analyzer_converter_last) begin
			main_rtio_analyzer_converter_mux <= 1'd0;
		end else begin
			main_rtio_analyzer_converter_mux <= (main_rtio_analyzer_converter_mux + 1'd1);
		end
	end
	if (main_rtio_analyzer_dma_reset_re) begin
		main_genericstandalone_interface1_bus_adr <= main_rtio_analyzer_dma_base_address_storage;
	end
	if (main_genericstandalone_interface1_bus_ack) begin
		if ((main_genericstandalone_interface1_bus_adr == main_rtio_analyzer_dma_last_address_storage)) begin
			main_genericstandalone_interface1_bus_adr <= main_rtio_analyzer_dma_base_address_storage;
		end else begin
			main_genericstandalone_interface1_bus_adr <= (main_genericstandalone_interface1_bus_adr + 1'd1);
		end
	end
	if (main_rtio_analyzer_dma_reset_re) begin
		main_rtio_analyzer_dma_message_count <= 1'd0;
	end
	if (main_genericstandalone_interface1_bus_ack) begin
		main_rtio_analyzer_dma_message_count <= (main_rtio_analyzer_dma_message_count + main_rtio_analyzer_dma_sink_payload_valid_token_count);
	end
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_cpulevel_arbiter_request[0])) begin
				if (builder_sdram_cpulevel_arbiter_request[1]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_cpulevel_arbiter_request[1])) begin
				if (builder_sdram_cpulevel_arbiter_request[0]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd0;
				end
			end
		end
	endcase
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_native_arbiter_request[0])) begin
				if (builder_sdram_native_arbiter_request[1]) begin
					builder_sdram_native_arbiter_grant <= 1'd1;
				end else begin
					if (builder_sdram_native_arbiter_request[2]) begin
						builder_sdram_native_arbiter_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_native_arbiter_request[1])) begin
				if (builder_sdram_native_arbiter_request[2]) begin
					builder_sdram_native_arbiter_grant <= 2'd2;
				end else begin
					if (builder_sdram_native_arbiter_request[0]) begin
						builder_sdram_native_arbiter_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~builder_sdram_native_arbiter_request[2])) begin
				if (builder_sdram_native_arbiter_request[0]) begin
					builder_sdram_native_arbiter_grant <= 1'd0;
				end else begin
					if (builder_sdram_native_arbiter_request[1]) begin
						builder_sdram_native_arbiter_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	case (builder_genericstandalone_grant)
		1'd0: begin
			if ((~builder_genericstandalone_request[0])) begin
				if (builder_genericstandalone_request[1]) begin
					builder_genericstandalone_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_genericstandalone_request[1])) begin
				if (builder_genericstandalone_request[0]) begin
					builder_genericstandalone_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_genericstandalone_slave_sel_r <= builder_genericstandalone_slave_sel;
	builder_genericstandalone_interface0_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank0_sel) begin
		case (builder_genericstandalone_interface0_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= builder_genericstandalone_csrbank0_dly_sel0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_w;
			end
			2'd2: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_w;
			end
			2'd3: begin
				builder_genericstandalone_interface0_bank_bus_dat_r <= main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank0_dly_sel0_re) begin
		main_genericstandalone_genericstandalone_ddrphy_storage_full[1:0] <= builder_genericstandalone_csrbank0_dly_sel0_r;
	end
	main_genericstandalone_genericstandalone_ddrphy_re <= builder_genericstandalone_csrbank0_dly_sel0_re;
	builder_genericstandalone_interface1_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank1_sel) begin
		case (builder_genericstandalone_interface1_bank_bus_adr[5:0])
			1'd0: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_control0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_command0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_address1_w;
			end
			3'd4: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_address0_w;
			end
			3'd5: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_baddress0_w;
			end
			3'd6: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_wrdata3_w;
			end
			3'd7: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_wrdata2_w;
			end
			4'd8: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_wrdata1_w;
			end
			4'd9: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_wrdata0_w;
			end
			4'd10: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_rddata3_w;
			end
			4'd11: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_rddata2_w;
			end
			4'd12: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_rddata1_w;
			end
			4'd13: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi0_rddata0_w;
			end
			4'd14: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_command0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_address1_w;
			end
			5'd17: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_address0_w;
			end
			5'd18: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_baddress0_w;
			end
			5'd19: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_wrdata3_w;
			end
			5'd20: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_wrdata2_w;
			end
			5'd21: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_wrdata1_w;
			end
			5'd22: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_wrdata0_w;
			end
			5'd23: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_rddata3_w;
			end
			5'd24: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_rddata2_w;
			end
			5'd25: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_rddata1_w;
			end
			5'd26: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi1_rddata0_w;
			end
			5'd27: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_command0_w;
			end
			5'd28: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_address1_w;
			end
			5'd30: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_address0_w;
			end
			5'd31: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_baddress0_w;
			end
			6'd32: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_wrdata3_w;
			end
			6'd33: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_wrdata2_w;
			end
			6'd34: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_wrdata1_w;
			end
			6'd35: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_wrdata0_w;
			end
			6'd36: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_rddata3_w;
			end
			6'd37: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_rddata2_w;
			end
			6'd38: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_rddata1_w;
			end
			6'd39: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi2_rddata0_w;
			end
			6'd40: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_command0_w;
			end
			6'd41: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_address1_w;
			end
			6'd43: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_address0_w;
			end
			6'd44: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_baddress0_w;
			end
			6'd45: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_wrdata3_w;
			end
			6'd46: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_wrdata2_w;
			end
			6'd47: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_wrdata1_w;
			end
			6'd48: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_wrdata0_w;
			end
			6'd49: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_rddata3_w;
			end
			6'd50: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_rddata2_w;
			end
			6'd51: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_rddata1_w;
			end
			6'd52: begin
				builder_genericstandalone_interface1_bank_bus_dat_r <= builder_genericstandalone_csrbank1_pi3_rddata0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank1_control0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_storage_full[3:0] <= builder_genericstandalone_csrbank1_control0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_re <= builder_genericstandalone_csrbank1_control0_re;
	if (builder_genericstandalone_csrbank1_pi0_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full[5:0] <= builder_genericstandalone_csrbank1_pi0_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re <= builder_genericstandalone_csrbank1_pi0_command0_re;
	if (builder_genericstandalone_csrbank1_pi0_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[14:8] <= builder_genericstandalone_csrbank1_pi0_address1_r;
	end
	if (builder_genericstandalone_csrbank1_pi0_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi0_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re <= builder_genericstandalone_csrbank1_pi0_address0_re;
	if (builder_genericstandalone_csrbank1_pi0_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank1_pi0_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re <= builder_genericstandalone_csrbank1_pi0_baddress0_re;
	if (builder_genericstandalone_csrbank1_pi0_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank1_pi0_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank1_pi0_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank1_pi0_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank1_pi0_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank1_pi0_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank1_pi0_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi0_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re <= builder_genericstandalone_csrbank1_pi0_wrdata0_re;
	if (builder_genericstandalone_csrbank1_pi1_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full[5:0] <= builder_genericstandalone_csrbank1_pi1_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re <= builder_genericstandalone_csrbank1_pi1_command0_re;
	if (builder_genericstandalone_csrbank1_pi1_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[14:8] <= builder_genericstandalone_csrbank1_pi1_address1_r;
	end
	if (builder_genericstandalone_csrbank1_pi1_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi1_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re <= builder_genericstandalone_csrbank1_pi1_address0_re;
	if (builder_genericstandalone_csrbank1_pi1_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank1_pi1_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re <= builder_genericstandalone_csrbank1_pi1_baddress0_re;
	if (builder_genericstandalone_csrbank1_pi1_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank1_pi1_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank1_pi1_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank1_pi1_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank1_pi1_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank1_pi1_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank1_pi1_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi1_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re <= builder_genericstandalone_csrbank1_pi1_wrdata0_re;
	if (builder_genericstandalone_csrbank1_pi2_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full[5:0] <= builder_genericstandalone_csrbank1_pi2_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re <= builder_genericstandalone_csrbank1_pi2_command0_re;
	if (builder_genericstandalone_csrbank1_pi2_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[14:8] <= builder_genericstandalone_csrbank1_pi2_address1_r;
	end
	if (builder_genericstandalone_csrbank1_pi2_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi2_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re <= builder_genericstandalone_csrbank1_pi2_address0_re;
	if (builder_genericstandalone_csrbank1_pi2_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank1_pi2_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re <= builder_genericstandalone_csrbank1_pi2_baddress0_re;
	if (builder_genericstandalone_csrbank1_pi2_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank1_pi2_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank1_pi2_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank1_pi2_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank1_pi2_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank1_pi2_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank1_pi2_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi2_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re <= builder_genericstandalone_csrbank1_pi2_wrdata0_re;
	if (builder_genericstandalone_csrbank1_pi3_command0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full[5:0] <= builder_genericstandalone_csrbank1_pi3_command0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re <= builder_genericstandalone_csrbank1_pi3_command0_re;
	if (builder_genericstandalone_csrbank1_pi3_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[14:8] <= builder_genericstandalone_csrbank1_pi3_address1_r;
	end
	if (builder_genericstandalone_csrbank1_pi3_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi3_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re <= builder_genericstandalone_csrbank1_pi3_address0_re;
	if (builder_genericstandalone_csrbank1_pi3_baddress0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full[2:0] <= builder_genericstandalone_csrbank1_pi3_baddress0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re <= builder_genericstandalone_csrbank1_pi3_baddress0_re;
	if (builder_genericstandalone_csrbank1_pi3_wrdata3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[31:24] <= builder_genericstandalone_csrbank1_pi3_wrdata3_r;
	end
	if (builder_genericstandalone_csrbank1_pi3_wrdata2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[23:16] <= builder_genericstandalone_csrbank1_pi3_wrdata2_r;
	end
	if (builder_genericstandalone_csrbank1_pi3_wrdata1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[15:8] <= builder_genericstandalone_csrbank1_pi3_wrdata1_r;
	end
	if (builder_genericstandalone_csrbank1_pi3_wrdata0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full[7:0] <= builder_genericstandalone_csrbank1_pi3_wrdata0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re <= builder_genericstandalone_csrbank1_pi3_wrdata0_re;
	builder_genericstandalone_interface2_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank2_sel) begin
		case (builder_genericstandalone_interface2_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_slot_w;
			end
			1'd1: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_length3_w;
			end
			2'd2: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_length2_w;
			end
			2'd3: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_length1_w;
			end
			3'd4: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_length0_w;
			end
			3'd5: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_errors3_w;
			end
			3'd6: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_errors2_w;
			end
			3'd7: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_errors1_w;
			end
			4'd8: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_errors0_w;
			end
			4'd9: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_writer_status_w;
			end
			4'd10: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_writer_pending_w;
			end
			4'd11: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_writer_ev_enable0_w;
			end
			4'd12: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_reader_start_w;
			end
			4'd13: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_reader_ready_w;
			end
			4'd14: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_reader_slot0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_reader_length1_w;
			end
			5'd16: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_reader_length0_w;
			end
			5'd17: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_reader_eventmanager_status_w;
			end
			5'd18: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= main_genericstandalone_reader_eventmanager_pending_w;
			end
			5'd19: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_sram_reader_ev_enable0_w;
			end
			5'd20: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_preamble_errors3_w;
			end
			5'd21: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_preamble_errors2_w;
			end
			5'd22: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_preamble_errors1_w;
			end
			5'd23: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_preamble_errors0_w;
			end
			5'd24: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_crc_errors3_w;
			end
			5'd25: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_crc_errors2_w;
			end
			5'd26: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_crc_errors1_w;
			end
			5'd27: begin
				builder_genericstandalone_interface2_bank_bus_dat_r <= builder_genericstandalone_csrbank2_crc_errors0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank2_sram_writer_ev_enable0_re) begin
		main_genericstandalone_writer_storage_full <= builder_genericstandalone_csrbank2_sram_writer_ev_enable0_r;
	end
	main_genericstandalone_writer_re <= builder_genericstandalone_csrbank2_sram_writer_ev_enable0_re;
	if (builder_genericstandalone_csrbank2_sram_reader_slot0_re) begin
		main_genericstandalone_reader_slot_storage_full[1:0] <= builder_genericstandalone_csrbank2_sram_reader_slot0_r;
	end
	main_genericstandalone_reader_slot_re <= builder_genericstandalone_csrbank2_sram_reader_slot0_re;
	if (builder_genericstandalone_csrbank2_sram_reader_length1_re) begin
		main_genericstandalone_reader_length_storage_full[10:8] <= builder_genericstandalone_csrbank2_sram_reader_length1_r;
	end
	if (builder_genericstandalone_csrbank2_sram_reader_length0_re) begin
		main_genericstandalone_reader_length_storage_full[7:0] <= builder_genericstandalone_csrbank2_sram_reader_length0_r;
	end
	main_genericstandalone_reader_length_re <= builder_genericstandalone_csrbank2_sram_reader_length0_re;
	if (builder_genericstandalone_csrbank2_sram_reader_ev_enable0_re) begin
		main_genericstandalone_reader_eventmanager_storage_full <= builder_genericstandalone_csrbank2_sram_reader_ev_enable0_r;
	end
	main_genericstandalone_reader_eventmanager_re <= builder_genericstandalone_csrbank2_sram_reader_ev_enable0_re;
	builder_genericstandalone_interface3_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank3_sel) begin
		case (builder_genericstandalone_interface3_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface3_bank_bus_dat_r <= builder_genericstandalone_csrbank3_in_w;
			end
			1'd1: begin
				builder_genericstandalone_interface3_bank_bus_dat_r <= builder_genericstandalone_csrbank3_out0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface3_bank_bus_dat_r <= builder_genericstandalone_csrbank3_oe0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank3_out0_re) begin
		main_i2c_out_storage_full[1:0] <= builder_genericstandalone_csrbank3_out0_r;
	end
	main_i2c_out_re <= builder_genericstandalone_csrbank3_out0_re;
	if (builder_genericstandalone_csrbank3_oe0_re) begin
		main_i2c_oe_storage_full[1:0] <= builder_genericstandalone_csrbank3_oe0_r;
	end
	main_i2c_oe_re <= builder_genericstandalone_csrbank3_oe0_re;
	builder_genericstandalone_interface4_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank4_sel) begin
		case (builder_genericstandalone_interface4_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_address0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface4_bank_bus_dat_r <= builder_genericstandalone_csrbank4_data_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank4_address0_re) begin
		main_add_identifier_storage_full[7:0] <= builder_genericstandalone_csrbank4_address0_r;
	end
	main_add_identifier_re <= builder_genericstandalone_csrbank4_address0_re;
	builder_genericstandalone_interface5_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank5_sel) begin
		case (builder_genericstandalone_interface5_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface5_bank_bus_dat_r <= builder_genericstandalone_csrbank5_reset0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank5_reset0_re) begin
		main_genericstandalone_kernel_cpu_storage_full <= builder_genericstandalone_csrbank5_reset0_r;
	end
	main_genericstandalone_kernel_cpu_re <= builder_genericstandalone_csrbank5_reset0_re;
	builder_genericstandalone_interface6_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank6_sel) begin
		case (builder_genericstandalone_interface6_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface6_bank_bus_dat_r <= builder_genericstandalone_csrbank6_out0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank6_out0_re) begin
		main_leds_storage_full <= builder_genericstandalone_csrbank6_out0_r;
	end
	main_leds_re <= builder_genericstandalone_csrbank6_out0_re;
	builder_genericstandalone_interface7_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank7_sel) begin
		case (builder_genericstandalone_interface7_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_enable0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_busy_w;
			end
			2'd2: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_message_encoder_overflow_w;
			end
			2'd3: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= main_rtio_analyzer_message_encoder_overflow_reset_w;
			end
			3'd4: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= main_rtio_analyzer_dma_reset_w;
			end
			3'd5: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_base_address4_w;
			end
			3'd6: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_base_address3_w;
			end
			3'd7: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_base_address2_w;
			end
			4'd8: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_base_address1_w;
			end
			4'd9: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_base_address0_w;
			end
			4'd10: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_last_address4_w;
			end
			4'd11: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_last_address3_w;
			end
			4'd12: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_last_address2_w;
			end
			4'd13: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_last_address1_w;
			end
			4'd14: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_last_address0_w;
			end
			4'd15: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count7_w;
			end
			5'd16: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count6_w;
			end
			5'd17: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count5_w;
			end
			5'd18: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count4_w;
			end
			5'd19: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count3_w;
			end
			5'd20: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count2_w;
			end
			5'd21: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count1_w;
			end
			5'd22: begin
				builder_genericstandalone_interface7_bank_bus_dat_r <= builder_genericstandalone_csrbank7_dma_byte_count0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank7_enable0_re) begin
		main_rtio_analyzer_enable_storage_full <= builder_genericstandalone_csrbank7_enable0_r;
	end
	main_rtio_analyzer_enable_re <= builder_genericstandalone_csrbank7_enable0_re;
	if (builder_genericstandalone_csrbank7_dma_base_address4_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[33:32] <= builder_genericstandalone_csrbank7_dma_base_address4_r;
	end
	if (builder_genericstandalone_csrbank7_dma_base_address3_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[31:24] <= builder_genericstandalone_csrbank7_dma_base_address3_r;
	end
	if (builder_genericstandalone_csrbank7_dma_base_address2_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[23:16] <= builder_genericstandalone_csrbank7_dma_base_address2_r;
	end
	if (builder_genericstandalone_csrbank7_dma_base_address1_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[15:8] <= builder_genericstandalone_csrbank7_dma_base_address1_r;
	end
	if (builder_genericstandalone_csrbank7_dma_base_address0_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[7:0] <= builder_genericstandalone_csrbank7_dma_base_address0_r;
	end
	main_rtio_analyzer_dma_base_address_re <= builder_genericstandalone_csrbank7_dma_base_address0_re;
	if (builder_genericstandalone_csrbank7_dma_last_address4_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[33:32] <= builder_genericstandalone_csrbank7_dma_last_address4_r;
	end
	if (builder_genericstandalone_csrbank7_dma_last_address3_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[31:24] <= builder_genericstandalone_csrbank7_dma_last_address3_r;
	end
	if (builder_genericstandalone_csrbank7_dma_last_address2_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[23:16] <= builder_genericstandalone_csrbank7_dma_last_address2_r;
	end
	if (builder_genericstandalone_csrbank7_dma_last_address1_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[15:8] <= builder_genericstandalone_csrbank7_dma_last_address1_r;
	end
	if (builder_genericstandalone_csrbank7_dma_last_address0_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[7:0] <= builder_genericstandalone_csrbank7_dma_last_address0_r;
	end
	main_rtio_analyzer_dma_last_address_re <= builder_genericstandalone_csrbank7_dma_last_address0_re;
	builder_genericstandalone_interface8_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank8_sel) begin
		case (builder_genericstandalone_interface8_bank_bus_adr[3:0])
			1'd0: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= main_rtio_core_reset_w;
			end
			1'd1: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= main_rtio_core_reset_phy_w;
			end
			2'd2: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= main_rtio_core_async_error_w;
			end
			2'd3: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_collision_channel1_w;
			end
			3'd4: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_collision_channel0_w;
			end
			3'd5: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_busy_channel1_w;
			end
			3'd6: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_busy_channel0_w;
			end
			3'd7: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_sequence_error_channel1_w;
			end
			4'd8: begin
				builder_genericstandalone_interface8_bank_bus_dat_r <= builder_genericstandalone_csrbank8_sequence_error_channel0_w;
			end
		endcase
	end
	builder_genericstandalone_interface9_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank9_sel) begin
		case (builder_genericstandalone_interface9_bank_bus_adr[0])
			1'd0: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_pll_reset0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface9_bank_bus_dat_r <= builder_genericstandalone_csrbank9_pll_locked_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank9_pll_reset0_re) begin
		main_rtio_crg_storage_full <= builder_genericstandalone_csrbank9_pll_reset0_r;
	end
	main_rtio_crg_re <= builder_genericstandalone_csrbank9_pll_reset0_re;
	builder_genericstandalone_interface10_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank10_sel) begin
		case (builder_genericstandalone_interface10_bank_bus_adr[2:0])
			1'd0: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_mon_chan_sel0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_mon_probe_sel0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= main_mon_value_update_w;
			end
			2'd3: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_mon_value_w;
			end
			3'd4: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_inj_chan_sel0_w;
			end
			3'd5: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= builder_genericstandalone_csrbank10_inj_override_sel0_w;
			end
			3'd6: begin
				builder_genericstandalone_interface10_bank_bus_dat_r <= main_inj_value_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank10_mon_chan_sel0_re) begin
		main_mon_chan_sel_storage_full[5:0] <= builder_genericstandalone_csrbank10_mon_chan_sel0_r;
	end
	main_mon_chan_sel_re <= builder_genericstandalone_csrbank10_mon_chan_sel0_re;
	if (builder_genericstandalone_csrbank10_mon_probe_sel0_re) begin
		main_mon_probe_sel_storage_full <= builder_genericstandalone_csrbank10_mon_probe_sel0_r;
	end
	main_mon_probe_sel_re <= builder_genericstandalone_csrbank10_mon_probe_sel0_re;
	if (builder_genericstandalone_csrbank10_inj_chan_sel0_re) begin
		main_inj_chan_sel_storage_full[5:0] <= builder_genericstandalone_csrbank10_inj_chan_sel0_r;
	end
	main_inj_chan_sel_re <= builder_genericstandalone_csrbank10_inj_chan_sel0_re;
	if (builder_genericstandalone_csrbank10_inj_override_sel0_re) begin
		main_inj_override_sel_storage_full[1:0] <= builder_genericstandalone_csrbank10_inj_override_sel0_r;
	end
	main_inj_override_sel_re <= builder_genericstandalone_csrbank10_inj_override_sel0_re;
	builder_genericstandalone_interface11_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank11_sel) begin
		case (builder_genericstandalone_interface11_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_bitbang0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_miso_w;
			end
			2'd2: begin
				builder_genericstandalone_interface11_bank_bus_dat_r <= builder_genericstandalone_csrbank11_bitbang_en0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank11_bitbang0_re) begin
		main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full[3:0] <= builder_genericstandalone_csrbank11_bitbang0_r;
	end
	main_genericstandalone_genericstandalone_spiflash_bitbang_re <= builder_genericstandalone_csrbank11_bitbang0_re;
	if (builder_genericstandalone_csrbank11_bitbang_en0_re) begin
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full <= builder_genericstandalone_csrbank11_bitbang_en0_r;
	end
	main_genericstandalone_genericstandalone_spiflash_bitbang_en_re <= builder_genericstandalone_csrbank11_bitbang_en0_re;
	builder_genericstandalone_interface12_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank12_sel) begin
		case (builder_genericstandalone_interface12_bank_bus_adr[4:0])
			1'd0: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load7_w;
			end
			1'd1: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load6_w;
			end
			2'd2: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load5_w;
			end
			2'd3: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load4_w;
			end
			3'd4: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load3_w;
			end
			3'd5: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load2_w;
			end
			3'd6: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load1_w;
			end
			3'd7: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_load0_w;
			end
			4'd8: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload7_w;
			end
			4'd9: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload6_w;
			end
			4'd10: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload5_w;
			end
			4'd11: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload4_w;
			end
			4'd12: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload3_w;
			end
			4'd13: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload2_w;
			end
			4'd14: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload1_w;
			end
			4'd15: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_reload0_w;
			end
			5'd16: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_en0_w;
			end
			5'd17: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_update_value_w;
			end
			5'd18: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value7_w;
			end
			5'd19: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value6_w;
			end
			5'd20: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value5_w;
			end
			5'd21: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value4_w;
			end
			5'd22: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value3_w;
			end
			5'd23: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value2_w;
			end
			5'd24: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value1_w;
			end
			5'd25: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_value0_w;
			end
			5'd26: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_status_w;
			end
			5'd27: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_pending_w;
			end
			5'd28: begin
				builder_genericstandalone_interface12_bank_bus_dat_r <= builder_genericstandalone_csrbank12_ev_enable0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank12_load7_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[63:56] <= builder_genericstandalone_csrbank12_load7_r;
	end
	if (builder_genericstandalone_csrbank12_load6_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[55:48] <= builder_genericstandalone_csrbank12_load6_r;
	end
	if (builder_genericstandalone_csrbank12_load5_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[47:40] <= builder_genericstandalone_csrbank12_load5_r;
	end
	if (builder_genericstandalone_csrbank12_load4_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[39:32] <= builder_genericstandalone_csrbank12_load4_r;
	end
	if (builder_genericstandalone_csrbank12_load3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[31:24] <= builder_genericstandalone_csrbank12_load3_r;
	end
	if (builder_genericstandalone_csrbank12_load2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[23:16] <= builder_genericstandalone_csrbank12_load2_r;
	end
	if (builder_genericstandalone_csrbank12_load1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[15:8] <= builder_genericstandalone_csrbank12_load1_r;
	end
	if (builder_genericstandalone_csrbank12_load0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full[7:0] <= builder_genericstandalone_csrbank12_load0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re <= builder_genericstandalone_csrbank12_load0_re;
	if (builder_genericstandalone_csrbank12_reload7_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[63:56] <= builder_genericstandalone_csrbank12_reload7_r;
	end
	if (builder_genericstandalone_csrbank12_reload6_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[55:48] <= builder_genericstandalone_csrbank12_reload6_r;
	end
	if (builder_genericstandalone_csrbank12_reload5_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[47:40] <= builder_genericstandalone_csrbank12_reload5_r;
	end
	if (builder_genericstandalone_csrbank12_reload4_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[39:32] <= builder_genericstandalone_csrbank12_reload4_r;
	end
	if (builder_genericstandalone_csrbank12_reload3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[31:24] <= builder_genericstandalone_csrbank12_reload3_r;
	end
	if (builder_genericstandalone_csrbank12_reload2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[23:16] <= builder_genericstandalone_csrbank12_reload2_r;
	end
	if (builder_genericstandalone_csrbank12_reload1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[15:8] <= builder_genericstandalone_csrbank12_reload1_r;
	end
	if (builder_genericstandalone_csrbank12_reload0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full[7:0] <= builder_genericstandalone_csrbank12_reload0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re <= builder_genericstandalone_csrbank12_reload0_re;
	if (builder_genericstandalone_csrbank12_en0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full <= builder_genericstandalone_csrbank12_en0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re <= builder_genericstandalone_csrbank12_en0_re;
	if (builder_genericstandalone_csrbank12_ev_enable0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full <= builder_genericstandalone_csrbank12_ev_enable0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re <= builder_genericstandalone_csrbank12_ev_enable0_re;
	builder_genericstandalone_interface13_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank13_sel) begin
		case (builder_genericstandalone_interface13_bank_bus_adr[2:0])
			1'd0: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_enable_null0_w;
			end
			1'd1: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_enable_prog0_w;
			end
			2'd2: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_prog_address3_w;
			end
			2'd3: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_prog_address2_w;
			end
			3'd4: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_prog_address1_w;
			end
			3'd5: begin
				builder_genericstandalone_interface13_bank_bus_dat_r <= builder_genericstandalone_csrbank13_prog_address0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank13_enable_null0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage_full <= builder_genericstandalone_csrbank13_enable_null0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_re <= builder_genericstandalone_csrbank13_enable_null0_re;
	if (builder_genericstandalone_csrbank13_enable_prog0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage_full <= builder_genericstandalone_csrbank13_enable_prog0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_re <= builder_genericstandalone_csrbank13_enable_prog0_re;
	if (builder_genericstandalone_csrbank13_prog_address3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[29:24] <= builder_genericstandalone_csrbank13_prog_address3_r;
	end
	if (builder_genericstandalone_csrbank13_prog_address2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[23:16] <= builder_genericstandalone_csrbank13_prog_address2_r;
	end
	if (builder_genericstandalone_csrbank13_prog_address1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[15:8] <= builder_genericstandalone_csrbank13_prog_address1_r;
	end
	if (builder_genericstandalone_csrbank13_prog_address0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full[7:0] <= builder_genericstandalone_csrbank13_prog_address0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_re <= builder_genericstandalone_csrbank13_prog_address0_re;
	builder_genericstandalone_interface14_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank14_sel) begin
		case (builder_genericstandalone_interface14_bank_bus_adr[2:0])
			1'd0: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_rxtx_w;
			end
			1'd1: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_txfull_w;
			end
			2'd2: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_rxempty_w;
			end
			2'd3: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_status_w;
			end
			3'd4: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= main_genericstandalone_genericstandalone_genericstandalone_uart_pending_w;
			end
			3'd5: begin
				builder_genericstandalone_interface14_bank_bus_dat_r <= builder_genericstandalone_csrbank14_ev_enable0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank14_ev_enable0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full[1:0] <= builder_genericstandalone_csrbank14_ev_enable0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_re <= builder_genericstandalone_csrbank14_ev_enable0_re;
	builder_genericstandalone_interface15_bank_bus_dat_r <= 1'd0;
	if (builder_genericstandalone_csrbank15_sel) begin
		case (builder_genericstandalone_interface15_bank_bus_adr[1:0])
			1'd0: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word3_w;
			end
			1'd1: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word2_w;
			end
			2'd2: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word1_w;
			end
			2'd3: begin
				builder_genericstandalone_interface15_bank_bus_dat_r <= builder_genericstandalone_csrbank15_tuning_word0_w;
			end
		endcase
	end
	if (builder_genericstandalone_csrbank15_tuning_word3_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[31:24] <= builder_genericstandalone_csrbank15_tuning_word3_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word2_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[23:16] <= builder_genericstandalone_csrbank15_tuning_word2_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word1_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[15:8] <= builder_genericstandalone_csrbank15_tuning_word1_r;
	end
	if (builder_genericstandalone_csrbank15_tuning_word0_re) begin
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full[7:0] <= builder_genericstandalone_csrbank15_tuning_word0_r;
	end
	main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re <= builder_genericstandalone_csrbank15_tuning_word0_re;
	if (sys_rst) begin
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_null_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_enable_prog_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_storage_full <= 30'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_prog_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_tmpu_error <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sram_bus_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_adr <= 14'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_we <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_interface_dat_w <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_dat_r <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_bus_wishbone_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_counter <= 2'd0;
		serial_tx <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_storage_full <= 32'd4367715;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_sink_ack <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_txen <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_tx <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_reg <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_bitcount <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_tx_busy <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_stb <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_source_payload_data <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_uart_clk_rxen <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_phase_accumulator_rx <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_r <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_reg <= 8'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_bitcount <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_phy_rx_busy <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_storage_full <= 2'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_level <= 5'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_produce <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_consume <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_level <= 5'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_produce <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_consume <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_storage_full <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_load_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_storage_full <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_reload_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_en_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value_status <= 64'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_pending <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_zero_old_trigger <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_eventmanager_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_timer0_value <= 64'd0;
		main_genericstandalone_genericstandalone_ddrphy_storage_full <= 2'd0;
		main_genericstandalone_genericstandalone_ddrphy_re <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_oe_dqs <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_oe_dq <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en0 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en1 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en2 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en3 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_n_rddata_en4 <= 1'd0;
		main_genericstandalone_genericstandalone_ddrphy_last_wrdata_en <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_storage_full <= 4'd0;
		main_genericstandalone_genericstandalone_genericstandalone_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector0_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector1_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector2_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_storage_full <= 6'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_command_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_storage_full <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_address_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_storage_full <= 3'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_baddress_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_storage_full <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_wrdata_re <= 1'd0;
		main_genericstandalone_genericstandalone_genericstandalone_phaseinjector3_status <= 32'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank0_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank1_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank2_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank3_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank4_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank5_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank6_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_idle <= 1'd1;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_bank7_row1 <= 15'd0;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_write2precharge_timer_count <= 3'd4;
		main_genericstandalone_genericstandalone_genericstandalone_sdram_controller_refresh_timer_count <= 10'd886;
		main_genericstandalone_genericstandalone_genericstandalone_adr_offset_r <= 2'd0;
		main_genericstandalone_genericstandalone_spiflash_bus_ack <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_storage_full <= 4'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_re <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_storage_full <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_bitbang_en_re <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_cs_n <= 1'd1;
		main_genericstandalone_genericstandalone_spiflash_clk <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_dq_oe <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_sr <= 32'd0;
		main_genericstandalone_genericstandalone_spiflash_i1 <= 1'd0;
		main_genericstandalone_genericstandalone_spiflash_dqi <= 2'd0;
		main_genericstandalone_genericstandalone_spiflash_counter <= 7'd0;
		main_genericstandalone_tx_mmcm_reset <= 1'd1;
		main_genericstandalone_rx_mmcm_reset <= 1'd1;
		main_genericstandalone_tx_init_qpll_reset0 <= 1'd0;
		main_genericstandalone_tx_init_tx_reset0 <= 1'd0;
		main_genericstandalone_tx_init_timer <= 6'd0;
		main_genericstandalone_tx_init_tick <= 1'd0;
		main_genericstandalone_rx_init_rx_reset0 <= 1'd0;
		main_genericstandalone_rx_init_drpvalue <= 16'd0;
		main_genericstandalone_rx_init_rx_pma_reset_done_r <= 1'd0;
		main_genericstandalone_cdr_lock_counter <= 13'd0;
		main_genericstandalone_cdr_locked <= 1'd0;
		main_genericstandalone_preamble_errors_status <= 32'd0;
		main_genericstandalone_crc_errors_status <= 32'd0;
		main_genericstandalone_tx_cdc_graycounter0_q <= 7'd0;
		main_genericstandalone_tx_cdc_graycounter0_q_binary <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter1_q <= 7'd0;
		main_genericstandalone_rx_cdc_graycounter1_q_binary <= 7'd0;
		main_genericstandalone_writer_errors_status <= 32'd0;
		main_genericstandalone_writer_storage_full <= 1'd0;
		main_genericstandalone_writer_re <= 1'd0;
		main_genericstandalone_writer_counter <= 32'd0;
		main_genericstandalone_writer_slot <= 2'd0;
		main_genericstandalone_writer_fifo_level <= 3'd0;
		main_genericstandalone_writer_fifo_produce <= 2'd0;
		main_genericstandalone_writer_fifo_consume <= 2'd0;
		main_genericstandalone_reader_slot_storage_full <= 2'd0;
		main_genericstandalone_reader_slot_re <= 1'd0;
		main_genericstandalone_reader_length_storage_full <= 11'd0;
		main_genericstandalone_reader_length_re <= 1'd0;
		main_genericstandalone_reader_done_pending <= 1'd0;
		main_genericstandalone_reader_eventmanager_storage_full <= 1'd0;
		main_genericstandalone_reader_eventmanager_re <= 1'd0;
		main_genericstandalone_reader_fifo_level <= 3'd0;
		main_genericstandalone_reader_fifo_produce <= 2'd0;
		main_genericstandalone_reader_fifo_consume <= 2'd0;
		main_genericstandalone_reader_counter <= 11'd0;
		main_genericstandalone_reader_last_d <= 1'd0;
		main_genericstandalone_sram0_bus_ack0 <= 1'd0;
		main_genericstandalone_sram1_bus_ack0 <= 1'd0;
		main_genericstandalone_sram2_bus_ack0 <= 1'd0;
		main_genericstandalone_sram3_bus_ack0 <= 1'd0;
		main_genericstandalone_sram0_bus_ack1 <= 1'd0;
		main_genericstandalone_sram1_bus_ack1 <= 1'd0;
		main_genericstandalone_sram2_bus_ack1 <= 1'd0;
		main_genericstandalone_sram3_bus_ack1 <= 1'd0;
		main_genericstandalone_slave_sel_r <= 8'd0;
		main_genericstandalone_kernel_cpu_storage_full <= 1'd1;
		main_genericstandalone_kernel_cpu_re <= 1'd0;
		main_genericstandalone_mailbox_i1_dat_r <= 32'd0;
		main_genericstandalone_mailbox_i1_ack <= 1'd0;
		main_genericstandalone_mailbox_i2_dat_r <= 32'd0;
		main_genericstandalone_mailbox_i2_ack <= 1'd0;
		main_genericstandalone_mailbox0 <= 32'd0;
		main_genericstandalone_mailbox1 <= 32'd0;
		main_genericstandalone_mailbox2 <= 32'd0;
		main_add_identifier_storage_full <= 8'd0;
		main_add_identifier_re <= 1'd0;
		main_leds_storage_full <= 1'd0;
		main_leds_re <= 1'd0;
		main_i2c_out_storage_full <= 2'd0;
		main_i2c_out_re <= 1'd0;
		main_i2c_oe_storage_full <= 2'd0;
		main_i2c_oe_re <= 1'd0;
		main_rtio_crg_storage_full <= 1'd1;
		main_rtio_crg_re <= 1'd0;
		main_rtio_core_collision_channel_status <= 16'd0;
		main_rtio_core_busy_channel_status <= 16'd0;
		main_rtio_core_sequence_error_channel_status <= 16'd0;
		main_rtio_core_cmd_reset <= 1'd1;
		main_rtio_core_cmd_reset_phy <= 1'd1;
		main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= 61'd0;
		main_rtio_core_o_collision <= 1'd0;
		main_rtio_core_o_busy <= 1'd0;
		main_rtio_core_o_sequence_error <= 1'd0;
		main_rtio_target_storage_full <= 32'd0;
		main_rtio_target_re <= 1'd0;
		main_rtio_o_data_storage_full <= 512'd0;
		main_rtio_o_data_re <= 1'd0;
		main_rtio_i_timeout_storage_full <= 64'd0;
		main_rtio_i_timeout_re <= 1'd0;
		main_rtio_counter_status <= 64'd0;
		main_rtio_now_hi_backing <= 32'd0;
		main_dma_dma_storage_full <= 34'd0;
		main_dma_dma_re <= 1'd0;
		main_dma_time_offset_storage_full <= 64'd0;
		main_dma_time_offset_re <= 1'd0;
		main_genericstandalone_csrbank0_bus_dat_r <= 32'd0;
		main_genericstandalone_csrbank0_bus_ack <= 1'd0;
		main_genericstandalone_csrbank1_bus_dat_r <= 32'd0;
		main_genericstandalone_csrbank1_bus_ack <= 1'd0;
		main_cri_con_storage_full <= 2'd0;
		main_cri_con_re <= 1'd0;
		main_cri_con_selected <= 1'd0;
		main_genericstandalone_csrbank2_bus_dat_r <= 32'd0;
		main_genericstandalone_csrbank2_bus_ack <= 1'd0;
		main_mon_chan_sel_storage_full <= 6'd0;
		main_mon_chan_sel_re <= 1'd0;
		main_mon_probe_sel_storage_full <= 1'd0;
		main_mon_probe_sel_re <= 1'd0;
		main_mon_status <= 1'd0;
		main_inj_chan_sel_storage_full <= 6'd0;
		main_inj_chan_sel_re <= 1'd0;
		main_inj_override_sel_storage_full <= 2'd0;
		main_inj_override_sel_re <= 1'd0;
		main_inj_o_sys0 <= 1'd0;
		main_inj_o_sys1 <= 1'd0;
		main_inj_o_sys2 <= 1'd0;
		main_inj_o_sys3 <= 1'd0;
		main_inj_o_sys4 <= 1'd0;
		main_inj_o_sys5 <= 1'd0;
		main_inj_o_sys6 <= 1'd0;
		main_inj_o_sys7 <= 1'd0;
		main_inj_o_sys8 <= 1'd0;
		main_inj_o_sys9 <= 1'd0;
		main_inj_o_sys10 <= 1'd0;
		main_inj_o_sys11 <= 1'd0;
		main_inj_o_sys12 <= 1'd0;
		main_inj_o_sys13 <= 1'd0;
		main_inj_o_sys14 <= 1'd0;
		main_inj_o_sys15 <= 1'd0;
		main_inj_o_sys16 <= 1'd0;
		main_inj_o_sys17 <= 1'd0;
		main_inj_o_sys18 <= 1'd0;
		main_inj_o_sys19 <= 1'd0;
		main_inj_o_sys20 <= 1'd0;
		main_inj_o_sys21 <= 1'd0;
		main_inj_o_sys22 <= 1'd0;
		main_inj_o_sys23 <= 1'd0;
		main_inj_o_sys24 <= 1'd0;
		main_inj_o_sys25 <= 1'd0;
		main_inj_o_sys26 <= 1'd0;
		main_inj_o_sys27 <= 1'd0;
		main_inj_o_sys28 <= 1'd0;
		main_inj_o_sys29 <= 1'd0;
		main_inj_o_sys30 <= 1'd0;
		main_inj_o_sys31 <= 1'd0;
		main_inj_o_sys32 <= 1'd0;
		main_inj_o_sys33 <= 1'd0;
		main_inj_o_sys34 <= 1'd0;
		main_inj_o_sys35 <= 1'd0;
		main_inj_o_sys36 <= 1'd0;
		main_inj_o_sys37 <= 1'd0;
		main_inj_o_sys38 <= 1'd0;
		main_inj_o_sys39 <= 1'd0;
		main_inj_o_sys40 <= 1'd0;
		main_inj_o_sys41 <= 1'd0;
		main_inj_o_sys42 <= 1'd0;
		main_inj_o_sys43 <= 1'd0;
		main_inj_o_sys44 <= 1'd0;
		main_inj_o_sys45 <= 1'd0;
		main_inj_o_sys46 <= 1'd0;
		main_inj_o_sys47 <= 1'd0;
		main_inj_o_sys48 <= 1'd0;
		main_inj_o_sys49 <= 1'd0;
		main_inj_o_sys50 <= 1'd0;
		main_inj_o_sys51 <= 1'd0;
		main_inj_o_sys52 <= 1'd0;
		main_inj_o_sys53 <= 1'd0;
		main_inj_o_sys54 <= 1'd0;
		main_inj_o_sys55 <= 1'd0;
		main_inj_o_sys56 <= 1'd0;
		main_inj_o_sys57 <= 1'd0;
		main_inj_o_sys58 <= 1'd0;
		main_inj_o_sys59 <= 1'd0;
		main_inj_o_sys60 <= 1'd0;
		main_inj_o_sys61 <= 1'd0;
		main_inj_o_sys62 <= 1'd0;
		main_inj_o_sys63 <= 1'd0;
		main_inj_o_sys64 <= 1'd0;
		main_inj_o_sys65 <= 1'd0;
		main_inj_o_sys66 <= 1'd0;
		main_inj_o_sys67 <= 1'd0;
		main_inj_o_sys68 <= 1'd0;
		main_inj_o_sys69 <= 1'd0;
		main_inj_o_sys70 <= 1'd0;
		main_inj_o_sys71 <= 1'd0;
		main_inj_o_sys72 <= 1'd0;
		main_inj_o_sys73 <= 1'd0;
		main_genericstandalone_interface1_bus_adr <= 30'd0;
		main_rtio_analyzer_enable_storage_full <= 1'd0;
		main_rtio_analyzer_enable_re <= 1'd0;
		main_rtio_analyzer_busy_status <= 1'd0;
		main_rtio_analyzer_message_encoder_source_stb <= 1'd0;
		main_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_rtio_analyzer_message_encoder_source_payload_data <= 256'd0;
		main_rtio_analyzer_message_encoder_status <= 1'd0;
		main_rtio_analyzer_message_encoder_read_wait_event_r <= 1'd0;
		main_rtio_analyzer_message_encoder_just_written <= 1'd0;
		main_rtio_analyzer_message_encoder_enable_r <= 1'd0;
		main_rtio_analyzer_message_encoder_stopping <= 1'd0;
		main_rtio_analyzer_fifo_readable <= 1'd0;
		main_rtio_analyzer_fifo_level0 <= 8'd0;
		main_rtio_analyzer_fifo_produce <= 7'd0;
		main_rtio_analyzer_fifo_consume <= 7'd0;
		main_rtio_analyzer_converter_mux <= 1'd0;
		main_rtio_analyzer_dma_base_address_storage_full <= 34'd0;
		main_rtio_analyzer_dma_base_address_re <= 1'd0;
		main_rtio_analyzer_dma_last_address_storage_full <= 34'd0;
		main_rtio_analyzer_dma_last_address_re <= 1'd0;
		main_rtio_analyzer_dma_message_count <= 59'd0;
		main_rtio_analyzer_enable_r <= 1'd0;
		builder_minicon_state <= 6'd0;
		builder_fullmemorywe_state <= 3'd0;
		builder_a7_1000basex_gtptxinit_state <= 2'd0;
		builder_a7_1000basex_gtprxinit_state <= 4'd0;
		builder_liteethmacsramwriter_state <= 2'd0;
		builder_liteethmacsramreader_state <= 2'd0;
		builder_grant <= 1'd0;
		builder_slave_sel_r <= 5'd0;
		builder_sdram_cpulevel_arbiter_grant <= 1'd0;
		builder_sdram_native_arbiter_grant <= 2'd0;
		builder_genericstandalone_grant <= 1'd0;
		builder_genericstandalone_slave_sel_r <= 6'd0;
		builder_genericstandalone_interface0_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface1_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface2_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface3_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface4_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface5_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface6_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface7_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface8_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface9_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface10_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface11_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface12_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface13_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface14_bank_bus_dat_r <= 8'd0;
		builder_genericstandalone_interface15_bank_bus_dat_r <= 8'd0;
	end
	builder_xilinxmultiregimpl0_regs0 <= serial_rx;
	builder_xilinxmultiregimpl0_regs1 <= builder_xilinxmultiregimpl0_regs0;
	builder_xilinxmultiregimpl4_regs0 <= main_genericstandalone_tx_init_qpll_lock0;
	builder_xilinxmultiregimpl4_regs1 <= builder_xilinxmultiregimpl4_regs0;
	builder_xilinxmultiregimpl5_regs0 <= main_genericstandalone_rx_init_rx_pma_reset_done0;
	builder_xilinxmultiregimpl5_regs1 <= builder_xilinxmultiregimpl5_regs0;
	builder_xilinxmultiregimpl6_regs0 <= main_genericstandalone_toggle_i;
	builder_xilinxmultiregimpl6_regs1 <= builder_xilinxmultiregimpl6_regs0;
	builder_xilinxmultiregimpl7_regs0 <= main_genericstandalone_ps_preamble_error_toggle_i;
	builder_xilinxmultiregimpl7_regs1 <= builder_xilinxmultiregimpl7_regs0;
	builder_xilinxmultiregimpl8_regs0 <= main_genericstandalone_ps_crc_error_toggle_i;
	builder_xilinxmultiregimpl8_regs1 <= builder_xilinxmultiregimpl8_regs0;
	builder_xilinxmultiregimpl10_regs0 <= main_genericstandalone_tx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl10_regs1 <= builder_xilinxmultiregimpl10_regs0;
	builder_xilinxmultiregimpl11_regs0 <= main_genericstandalone_rx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl11_regs1 <= builder_xilinxmultiregimpl11_regs0;
	builder_xilinxmultiregimpl13_regs0 <= main_i2c_tstriple0_i;
	builder_xilinxmultiregimpl13_regs1 <= builder_xilinxmultiregimpl13_regs0;
	builder_xilinxmultiregimpl14_regs0 <= main_i2c_tstriple1_i;
	builder_xilinxmultiregimpl14_regs1 <= builder_xilinxmultiregimpl14_regs0;
	builder_xilinxmultiregimpl15_regs0 <= main_rtio_crg_pll_locked;
	builder_xilinxmultiregimpl15_regs1 <= builder_xilinxmultiregimpl15_regs0;
	builder_xilinxmultiregimpl16_regs0 <= main_rtio_tsc_value_gray_rtio;
	builder_xilinxmultiregimpl16_regs1 <= builder_xilinxmultiregimpl16_regs0;
	builder_xilinxmultiregimpl83_regs0 <= main_mon_bussynchronizer0_i;
	builder_xilinxmultiregimpl83_regs1 <= builder_xilinxmultiregimpl83_regs0;
	builder_xilinxmultiregimpl84_regs0 <= main_mon_bussynchronizer1_i;
	builder_xilinxmultiregimpl84_regs1 <= builder_xilinxmultiregimpl84_regs0;
	builder_xilinxmultiregimpl85_regs0 <= main_mon_bussynchronizer2_i;
	builder_xilinxmultiregimpl85_regs1 <= builder_xilinxmultiregimpl85_regs0;
	builder_xilinxmultiregimpl86_regs0 <= main_mon_bussynchronizer3_i;
	builder_xilinxmultiregimpl86_regs1 <= builder_xilinxmultiregimpl86_regs0;
	builder_xilinxmultiregimpl87_regs0 <= main_mon_bussynchronizer4_i;
	builder_xilinxmultiregimpl87_regs1 <= builder_xilinxmultiregimpl87_regs0;
	builder_xilinxmultiregimpl88_regs0 <= main_mon_bussynchronizer5_i;
	builder_xilinxmultiregimpl88_regs1 <= builder_xilinxmultiregimpl88_regs0;
	builder_xilinxmultiregimpl89_regs0 <= main_mon_bussynchronizer6_i;
	builder_xilinxmultiregimpl89_regs1 <= builder_xilinxmultiregimpl89_regs0;
	builder_xilinxmultiregimpl90_regs0 <= main_mon_bussynchronizer7_i;
	builder_xilinxmultiregimpl90_regs1 <= builder_xilinxmultiregimpl90_regs0;
	builder_xilinxmultiregimpl91_regs0 <= main_mon_bussynchronizer8_i;
	builder_xilinxmultiregimpl91_regs1 <= builder_xilinxmultiregimpl91_regs0;
	builder_xilinxmultiregimpl92_regs0 <= main_mon_bussynchronizer9_i;
	builder_xilinxmultiregimpl92_regs1 <= builder_xilinxmultiregimpl92_regs0;
	builder_xilinxmultiregimpl93_regs0 <= main_mon_bussynchronizer10_i;
	builder_xilinxmultiregimpl93_regs1 <= builder_xilinxmultiregimpl93_regs0;
	builder_xilinxmultiregimpl94_regs0 <= main_mon_bussynchronizer11_i;
	builder_xilinxmultiregimpl94_regs1 <= builder_xilinxmultiregimpl94_regs0;
	builder_xilinxmultiregimpl95_regs0 <= main_mon_bussynchronizer12_i;
	builder_xilinxmultiregimpl95_regs1 <= builder_xilinxmultiregimpl95_regs0;
	builder_xilinxmultiregimpl96_regs0 <= main_mon_bussynchronizer13_i;
	builder_xilinxmultiregimpl96_regs1 <= builder_xilinxmultiregimpl96_regs0;
	builder_xilinxmultiregimpl97_regs0 <= main_mon_bussynchronizer14_i;
	builder_xilinxmultiregimpl97_regs1 <= builder_xilinxmultiregimpl97_regs0;
	builder_xilinxmultiregimpl98_regs0 <= main_mon_bussynchronizer15_i;
	builder_xilinxmultiregimpl98_regs1 <= builder_xilinxmultiregimpl98_regs0;
	builder_xilinxmultiregimpl99_regs0 <= main_mon_bussynchronizer16_i;
	builder_xilinxmultiregimpl99_regs1 <= builder_xilinxmultiregimpl99_regs0;
	builder_xilinxmultiregimpl100_regs0 <= main_mon_bussynchronizer17_i;
	builder_xilinxmultiregimpl100_regs1 <= builder_xilinxmultiregimpl100_regs0;
	builder_xilinxmultiregimpl101_regs0 <= main_mon_bussynchronizer18_i;
	builder_xilinxmultiregimpl101_regs1 <= builder_xilinxmultiregimpl101_regs0;
	builder_xilinxmultiregimpl102_regs0 <= main_mon_bussynchronizer19_i;
	builder_xilinxmultiregimpl102_regs1 <= builder_xilinxmultiregimpl102_regs0;
	builder_xilinxmultiregimpl103_regs0 <= main_mon_bussynchronizer20_i;
	builder_xilinxmultiregimpl103_regs1 <= builder_xilinxmultiregimpl103_regs0;
	builder_xilinxmultiregimpl104_regs0 <= main_mon_bussynchronizer21_i;
	builder_xilinxmultiregimpl104_regs1 <= builder_xilinxmultiregimpl104_regs0;
	builder_xilinxmultiregimpl105_regs0 <= main_mon_bussynchronizer22_i;
	builder_xilinxmultiregimpl105_regs1 <= builder_xilinxmultiregimpl105_regs0;
	builder_xilinxmultiregimpl106_regs0 <= main_mon_bussynchronizer23_i;
	builder_xilinxmultiregimpl106_regs1 <= builder_xilinxmultiregimpl106_regs0;
	builder_xilinxmultiregimpl107_regs0 <= main_mon_bussynchronizer24_i;
	builder_xilinxmultiregimpl107_regs1 <= builder_xilinxmultiregimpl107_regs0;
	builder_xilinxmultiregimpl108_regs0 <= main_mon_bussynchronizer25_i;
	builder_xilinxmultiregimpl108_regs1 <= builder_xilinxmultiregimpl108_regs0;
	builder_xilinxmultiregimpl109_regs0 <= main_mon_bussynchronizer26_i;
	builder_xilinxmultiregimpl109_regs1 <= builder_xilinxmultiregimpl109_regs0;
	builder_xilinxmultiregimpl110_regs0 <= main_mon_bussynchronizer27_i;
	builder_xilinxmultiregimpl110_regs1 <= builder_xilinxmultiregimpl110_regs0;
	builder_xilinxmultiregimpl111_regs0 <= main_mon_bussynchronizer28_i;
	builder_xilinxmultiregimpl111_regs1 <= builder_xilinxmultiregimpl111_regs0;
	builder_xilinxmultiregimpl112_regs0 <= main_mon_bussynchronizer29_i;
	builder_xilinxmultiregimpl112_regs1 <= builder_xilinxmultiregimpl112_regs0;
	builder_xilinxmultiregimpl113_regs0 <= main_mon_bussynchronizer30_i;
	builder_xilinxmultiregimpl113_regs1 <= builder_xilinxmultiregimpl113_regs0;
	builder_xilinxmultiregimpl114_regs0 <= main_mon_bussynchronizer31_i;
	builder_xilinxmultiregimpl114_regs1 <= builder_xilinxmultiregimpl114_regs0;
	builder_xilinxmultiregimpl115_regs0 <= main_mon_bussynchronizer32_i;
	builder_xilinxmultiregimpl115_regs1 <= builder_xilinxmultiregimpl115_regs0;
	builder_xilinxmultiregimpl116_regs0 <= main_mon_bussynchronizer33_i;
	builder_xilinxmultiregimpl116_regs1 <= builder_xilinxmultiregimpl116_regs0;
	builder_xilinxmultiregimpl117_regs0 <= main_mon_bussynchronizer34_i;
	builder_xilinxmultiregimpl117_regs1 <= builder_xilinxmultiregimpl117_regs0;
	builder_xilinxmultiregimpl118_regs0 <= main_mon_bussynchronizer35_i;
	builder_xilinxmultiregimpl118_regs1 <= builder_xilinxmultiregimpl118_regs0;
	builder_xilinxmultiregimpl119_regs0 <= main_mon_bussynchronizer36_i;
	builder_xilinxmultiregimpl119_regs1 <= builder_xilinxmultiregimpl119_regs0;
	builder_xilinxmultiregimpl120_regs0 <= main_mon_bussynchronizer37_i;
	builder_xilinxmultiregimpl120_regs1 <= builder_xilinxmultiregimpl120_regs0;
	builder_xilinxmultiregimpl121_regs0 <= main_mon_bussynchronizer38_i;
	builder_xilinxmultiregimpl121_regs1 <= builder_xilinxmultiregimpl121_regs0;
	builder_xilinxmultiregimpl122_regs0 <= main_mon_bussynchronizer39_i;
	builder_xilinxmultiregimpl122_regs1 <= builder_xilinxmultiregimpl122_regs0;
	builder_xilinxmultiregimpl123_regs0 <= main_mon_bussynchronizer40_i;
	builder_xilinxmultiregimpl123_regs1 <= builder_xilinxmultiregimpl123_regs0;
end

always @(posedge sys_kernel_clk) begin
	main_dma_dma_enable_r <= main_dma_flow_enable;
	if ((main_dma_flow_enable & (~main_dma_dma_enable_r))) begin
		main_dma_dma_sink_payload_address <= main_dma_dma_storage;
		main_dma_dma_sink_eop <= 1'd0;
		main_dma_dma_sink_stb <= 1'd1;
	end
	if ((main_dma_dma_sink_stb & main_dma_dma_sink_ack)) begin
		if (main_dma_dma_sink_eop) begin
			main_dma_dma_sink_stb <= 1'd0;
		end else begin
			main_dma_dma_sink_payload_address <= (main_dma_dma_sink_payload_address + 1'd1);
			if ((~main_dma_flow_enable)) begin
				main_dma_dma_sink_eop <= 1'd1;
			end
		end
	end
	if (main_dma_dma_source_ack) begin
		main_dma_dma_data_reg_loaded <= 1'd0;
	end
	if (main_genericstandalone_interface0_bus_ack) begin
		main_dma_dma_data_reg_loaded <= 1'd1;
		main_dma_dma_source_payload_data <= main_genericstandalone_interface0_bus_dat_r;
		main_dma_dma_source_eop <= main_dma_dma_sink_eop;
	end
	main_dma_rawslicer_level <= main_dma_rawslicer_next_level;
	if (main_dma_rawslicer_load_buf) begin
		case (main_dma_rawslicer_level)
			1'd0: begin
				main_dma_rawslicer_buf[127:0] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			1'd1: begin
				main_dma_rawslicer_buf[135:8] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd2: begin
				main_dma_rawslicer_buf[143:16] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd3: begin
				main_dma_rawslicer_buf[151:24] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd4: begin
				main_dma_rawslicer_buf[159:32] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd5: begin
				main_dma_rawslicer_buf[167:40] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd6: begin
				main_dma_rawslicer_buf[175:48] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd7: begin
				main_dma_rawslicer_buf[183:56] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd8: begin
				main_dma_rawslicer_buf[191:64] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd9: begin
				main_dma_rawslicer_buf[199:72] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd10: begin
				main_dma_rawslicer_buf[207:80] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd11: begin
				main_dma_rawslicer_buf[215:88] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd12: begin
				main_dma_rawslicer_buf[223:96] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd13: begin
				main_dma_rawslicer_buf[231:104] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd14: begin
				main_dma_rawslicer_buf[239:112] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd15: begin
				main_dma_rawslicer_buf[247:120] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd16: begin
				main_dma_rawslicer_buf[255:128] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd17: begin
				main_dma_rawslicer_buf[263:136] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd18: begin
				main_dma_rawslicer_buf[271:144] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd19: begin
				main_dma_rawslicer_buf[279:152] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd20: begin
				main_dma_rawslicer_buf[287:160] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd21: begin
				main_dma_rawslicer_buf[295:168] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd22: begin
				main_dma_rawslicer_buf[303:176] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd23: begin
				main_dma_rawslicer_buf[311:184] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd24: begin
				main_dma_rawslicer_buf[319:192] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd25: begin
				main_dma_rawslicer_buf[327:200] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd26: begin
				main_dma_rawslicer_buf[335:208] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd27: begin
				main_dma_rawslicer_buf[343:216] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd28: begin
				main_dma_rawslicer_buf[351:224] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd29: begin
				main_dma_rawslicer_buf[359:232] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd30: begin
				main_dma_rawslicer_buf[367:240] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd31: begin
				main_dma_rawslicer_buf[375:248] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd32: begin
				main_dma_rawslicer_buf[383:256] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd33: begin
				main_dma_rawslicer_buf[391:264] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd34: begin
				main_dma_rawslicer_buf[399:272] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd35: begin
				main_dma_rawslicer_buf[407:280] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd36: begin
				main_dma_rawslicer_buf[415:288] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd37: begin
				main_dma_rawslicer_buf[423:296] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd38: begin
				main_dma_rawslicer_buf[431:304] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd39: begin
				main_dma_rawslicer_buf[439:312] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd40: begin
				main_dma_rawslicer_buf[447:320] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd41: begin
				main_dma_rawslicer_buf[455:328] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd42: begin
				main_dma_rawslicer_buf[463:336] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd43: begin
				main_dma_rawslicer_buf[471:344] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd44: begin
				main_dma_rawslicer_buf[479:352] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd45: begin
				main_dma_rawslicer_buf[487:360] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd46: begin
				main_dma_rawslicer_buf[495:368] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd47: begin
				main_dma_rawslicer_buf[503:376] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd48: begin
				main_dma_rawslicer_buf[511:384] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd49: begin
				main_dma_rawslicer_buf[519:392] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd50: begin
				main_dma_rawslicer_buf[527:400] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd51: begin
				main_dma_rawslicer_buf[535:408] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd52: begin
				main_dma_rawslicer_buf[543:416] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd53: begin
				main_dma_rawslicer_buf[551:424] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd54: begin
				main_dma_rawslicer_buf[559:432] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd55: begin
				main_dma_rawslicer_buf[567:440] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd56: begin
				main_dma_rawslicer_buf[575:448] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd57: begin
				main_dma_rawslicer_buf[583:456] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd58: begin
				main_dma_rawslicer_buf[591:464] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd59: begin
				main_dma_rawslicer_buf[599:472] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd60: begin
				main_dma_rawslicer_buf[607:480] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd61: begin
				main_dma_rawslicer_buf[615:488] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd62: begin
				main_dma_rawslicer_buf[623:496] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd63: begin
				main_dma_rawslicer_buf[631:504] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd64: begin
				main_dma_rawslicer_buf[639:512] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd65: begin
				main_dma_rawslicer_buf[647:520] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd66: begin
				main_dma_rawslicer_buf[655:528] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd67: begin
				main_dma_rawslicer_buf[663:536] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd68: begin
				main_dma_rawslicer_buf[671:544] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd69: begin
				main_dma_rawslicer_buf[679:552] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd70: begin
				main_dma_rawslicer_buf[687:560] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd71: begin
				main_dma_rawslicer_buf[695:568] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd72: begin
				main_dma_rawslicer_buf[703:576] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd73: begin
				main_dma_rawslicer_buf[711:584] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd74: begin
				main_dma_rawslicer_buf[719:592] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd75: begin
				main_dma_rawslicer_buf[727:600] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd76: begin
				main_dma_rawslicer_buf[735:608] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120]};
			end
		endcase
	end
	if (main_dma_rawslicer_shift_buf) begin
		case (main_dma_rawslicer_source_consume)
			1'd0: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:0];
			end
			1'd1: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:8];
			end
			2'd2: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:16];
			end
			2'd3: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:24];
			end
			3'd4: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:32];
			end
			3'd5: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:40];
			end
			3'd6: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:48];
			end
			3'd7: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:56];
			end
			4'd8: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:64];
			end
			4'd9: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:72];
			end
			4'd10: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:80];
			end
			4'd11: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:88];
			end
			4'd12: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:96];
			end
			4'd13: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:104];
			end
			4'd14: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:112];
			end
			4'd15: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:120];
			end
			5'd16: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:128];
			end
			5'd17: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:136];
			end
			5'd18: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:144];
			end
			5'd19: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:152];
			end
			5'd20: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:160];
			end
			5'd21: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:168];
			end
			5'd22: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:176];
			end
			5'd23: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:184];
			end
			5'd24: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:192];
			end
			5'd25: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:200];
			end
			5'd26: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:208];
			end
			5'd27: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:216];
			end
			5'd28: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:224];
			end
			5'd29: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:232];
			end
			5'd30: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:240];
			end
			5'd31: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:248];
			end
			6'd32: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:256];
			end
			6'd33: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:264];
			end
			6'd34: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:272];
			end
			6'd35: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:280];
			end
			6'd36: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:288];
			end
			6'd37: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:296];
			end
			6'd38: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:304];
			end
			6'd39: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:312];
			end
			6'd40: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:320];
			end
			6'd41: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:328];
			end
			6'd42: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:336];
			end
			6'd43: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:344];
			end
			6'd44: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:352];
			end
			6'd45: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:360];
			end
			6'd46: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:368];
			end
			6'd47: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:376];
			end
			6'd48: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:384];
			end
			6'd49: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:392];
			end
			6'd50: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:400];
			end
			6'd51: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:408];
			end
			6'd52: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:416];
			end
			6'd53: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:424];
			end
			6'd54: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:432];
			end
			6'd55: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:440];
			end
			6'd56: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:448];
			end
			6'd57: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:456];
			end
			6'd58: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:464];
			end
			6'd59: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:472];
			end
			6'd60: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:480];
			end
			6'd61: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:488];
			end
			6'd62: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:496];
			end
			6'd63: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:504];
			end
			7'd64: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:512];
			end
			7'd65: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:520];
			end
			7'd66: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:528];
			end
			7'd67: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:536];
			end
			7'd68: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:544];
			end
			7'd69: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:552];
			end
			7'd70: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:560];
			end
			7'd71: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:568];
			end
			7'd72: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:576];
			end
			7'd73: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:584];
			end
			7'd74: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:592];
			end
			7'd75: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:600];
			end
			7'd76: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[735:608];
			end
		endcase
	end
	builder_clockdomainsrenamer_resetinserter_state <= builder_clockdomainsrenamer_resetinserter_next_state;
	if (main_dma_reset) begin
		main_dma_rawslicer_buf <= 736'd0;
		main_dma_rawslicer_level <= 7'd0;
		builder_clockdomainsrenamer_resetinserter_state <= 2'd0;
	end
	builder_clockdomainsrenamer_recordconverter_state <= builder_clockdomainsrenamer_recordconverter_next_state;
	if (main_dma_time_offset_source_ack) begin
		main_dma_time_offset_source_stb <= 1'd0;
	end
	if ((~main_dma_time_offset_source_stb)) begin
		main_dma_time_offset_source_payload_length <= main_dma_time_offset_sink_payload_length;
		main_dma_time_offset_source_payload_channel <= main_dma_time_offset_sink_payload_channel;
		main_dma_time_offset_source_payload_address <= main_dma_time_offset_sink_payload_address;
		main_dma_time_offset_source_payload_data <= main_dma_time_offset_sink_payload_data;
		main_dma_time_offset_source_payload_timestamp <= (main_dma_time_offset_sink_payload_timestamp + main_dma_time_offset_storage);
		main_dma_time_offset_source_eop <= main_dma_time_offset_sink_eop;
		main_dma_time_offset_source_stb <= main_dma_time_offset_sink_stb;
	end
	if (main_dma_cri_master_underflow_trigger) begin
		main_dma_cri_master_error_w <= 1'd1;
		main_dma_cri_master_error_channel_status <= main_dma_cri_master_sink_payload_channel;
		main_dma_cri_master_error_timestamp_status <= main_dma_cri_master_sink_payload_timestamp;
		main_dma_cri_master_error_address_status <= main_dma_cri_master_sink_payload_address;
	end
	if (main_dma_cri_master_link_error_trigger) begin
		main_dma_cri_master_error_w <= 2'd2;
		main_dma_cri_master_error_channel_status <= main_dma_cri_master_sink_payload_channel;
		main_dma_cri_master_error_timestamp_status <= main_dma_cri_master_sink_payload_timestamp;
		main_dma_cri_master_error_address_status <= main_dma_cri_master_sink_payload_address;
	end
	if (main_dma_cri_master_error_re) begin
		main_dma_cri_master_error_w <= 1'd0;
	end
	builder_clockdomainsrenamer_crimaster_state <= builder_clockdomainsrenamer_crimaster_next_state;
	builder_clockdomainsrenamer_fsm_state <= builder_clockdomainsrenamer_fsm_next_state;
	if (sys_kernel_rst) begin
		main_dma_dma_sink_stb <= 1'd0;
		main_dma_dma_sink_eop <= 1'd0;
		main_dma_dma_sink_payload_address <= 30'd0;
		main_dma_dma_source_eop <= 1'd0;
		main_dma_dma_source_payload_data <= 128'd0;
		main_dma_dma_data_reg_loaded <= 1'd0;
		main_dma_dma_enable_r <= 1'd0;
		main_dma_rawslicer_buf <= 736'd0;
		main_dma_rawslicer_level <= 7'd0;
		main_dma_time_offset_source_stb <= 1'd0;
		main_dma_time_offset_source_eop <= 1'd0;
		main_dma_time_offset_source_payload_length <= 8'd0;
		main_dma_time_offset_source_payload_channel <= 24'd0;
		main_dma_time_offset_source_payload_timestamp <= 64'd0;
		main_dma_time_offset_source_payload_address <= 8'd0;
		main_dma_time_offset_source_payload_data <= 512'd0;
		main_dma_cri_master_error_w <= 2'd0;
		main_dma_cri_master_error_channel_status <= 24'd0;
		main_dma_cri_master_error_timestamp_status <= 64'd0;
		main_dma_cri_master_error_address_status <= 16'd0;
		builder_clockdomainsrenamer_resetinserter_state <= 2'd0;
		builder_clockdomainsrenamer_recordconverter_state <= 2'd0;
		builder_clockdomainsrenamer_crimaster_state <= 3'd0;
		builder_clockdomainsrenamer_fsm_state <= 3'd0;
	end
end

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(23'd4194304)
) mor1kx (
	.clk(sys_clk),
	.dwbm_ack_i(main_genericstandalone_genericstandalone_genericstandalone_dbus_ack),
	.dwbm_dat_i(main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_r),
	.dwbm_err_i(main_genericstandalone_genericstandalone_genericstandalone_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(main_genericstandalone_genericstandalone_genericstandalone_interrupt),
	.iwbm_ack_i(main_genericstandalone_genericstandalone_genericstandalone_ibus_ack),
	.iwbm_dat_i(main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_r),
	.iwbm_err_i(main_genericstandalone_genericstandalone_genericstandalone_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_rst),
	.dwbm_adr_o(main_genericstandalone_genericstandalone_genericstandalone_d_adr_o),
	.dwbm_bte_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_bte),
	.dwbm_cti_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_cti),
	.dwbm_cyc_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_cyc),
	.dwbm_dat_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_dat_w),
	.dwbm_sel_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_sel),
	.dwbm_stb_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_stb),
	.dwbm_we_o(main_genericstandalone_genericstandalone_genericstandalone_dbus_we),
	.iwbm_adr_o(main_genericstandalone_genericstandalone_genericstandalone_i_adr_o),
	.iwbm_bte_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_bte),
	.iwbm_cti_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_cti),
	.iwbm_cyc_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_cyc),
	.iwbm_dat_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_dat_w),
	.iwbm_sel_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_sel),
	.iwbm_stb_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_stb),
	.iwbm_we_o(main_genericstandalone_genericstandalone_genericstandalone_ibus_we)
);

reg [31:0] mem[0:1023];
reg [9:0] memadr;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_sram_we[0])
		mem[main_genericstandalone_genericstandalone_genericstandalone_sram_adr][7:0] <= main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w[7:0];
	if (main_genericstandalone_genericstandalone_genericstandalone_sram_we[1])
		mem[main_genericstandalone_genericstandalone_genericstandalone_sram_adr][15:8] <= main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w[15:8];
	if (main_genericstandalone_genericstandalone_genericstandalone_sram_we[2])
		mem[main_genericstandalone_genericstandalone_genericstandalone_sram_adr][23:16] <= main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w[23:16];
	if (main_genericstandalone_genericstandalone_genericstandalone_sram_we[3])
		mem[main_genericstandalone_genericstandalone_genericstandalone_sram_adr][31:24] <= main_genericstandalone_genericstandalone_genericstandalone_sram_dat_w[31:24];
	memadr <= main_genericstandalone_genericstandalone_genericstandalone_sram_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_sram_dat_r = mem[memadr];

reg [8:0] storage[0:15];
reg [8:0] memdat;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_we)
		storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr] <= main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_wrport_dat_r = memdat;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_dat_r = storage[main_genericstandalone_genericstandalone_genericstandalone_uart_tx_fifo_rdport_adr];

reg [8:0] storage_1[0:15];
reg [8:0] memdat_1;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_we)
		storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr] <= main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_w;
	memdat_1 <= storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_wrport_dat_r = memdat_1;
assign main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_dat_r = storage_1[main_genericstandalone_genericstandalone_genericstandalone_uart_rx_fifo_rdport_adr];

IBUFDS_GTE2 IBUFDS_GTE2(
	.CEB(1'd0),
	.I(clk125_gtp_p),
	.IB(clk125_gtp_n),
	.O(main_genericstandalone_genericstandalone_clk125_buf),
	.ODIV2(main_genericstandalone_genericstandalone_clk125_div2)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(14.5),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(8.0),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(90.0),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE (
	.CLKFBIN(main_genericstandalone_genericstandalone_mmcm_fb),
	.CLKIN1(main_genericstandalone_genericstandalone_clk125_div2),
	.CLKFBOUT(main_genericstandalone_genericstandalone_mmcm_fb),
	.CLKOUT0(main_genericstandalone_genericstandalone_mmcm_sys),
	.CLKOUT1(main_genericstandalone_genericstandalone_mmcm_sys4x),
	.CLKOUT2(main_genericstandalone_genericstandalone_mmcm_sys4x_dqs),
	.LOCKED(main_genericstandalone_genericstandalone_mmcm_locked)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE(3'd5),
	.CLKOUT0_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1)
) PLLE2_BASE (
	.CLKFBIN(main_genericstandalone_genericstandalone_pll_fb),
	.CLKIN1(main_genericstandalone_genericstandalone_clk125_div2),
	.CLKFBOUT(main_genericstandalone_genericstandalone_pll_fb),
	.CLKOUT0(main_genericstandalone_genericstandalone_pll_clk200),
	.LOCKED(main_genericstandalone_genericstandalone_pll_locked)
);

BUFG BUFG(
	.I(main_genericstandalone_genericstandalone_mmcm_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(main_genericstandalone_genericstandalone_mmcm_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_2(
	.I(main_genericstandalone_genericstandalone_mmcm_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

BUFG BUFG_3(
	.I(main_genericstandalone_genericstandalone_pll_clk200),
	.O(clk200_clk)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg),
	.Q(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_meta),
	.PRE(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg),
	.Q(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_unbuf)
);

BUFG BUFG_4(
	.I(main_genericstandalone_genericstandalone_asyncresetsynchronizerbufg_rst_unbuf),
	.O(sys_rst)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(main_genericstandalone_genericstandalone_ic_reset)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(main_genericstandalone_genericstandalone_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[0]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[0]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[0]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[1]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[1]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[3]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[3]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[3]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[3]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[3]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[3]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[4]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[4]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[4]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[4]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[4]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[4]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[5]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[5]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[5]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[5]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[5]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[5]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[6]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[6]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[6]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[6]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[6]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[6]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[7]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[7]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[7]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[7]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[7]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[7]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[7]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[8]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[8]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[8]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[8]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[8]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[8]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[8]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[9]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[9]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[9]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[9]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[9]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[9]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[9]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[10]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[10]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[10]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[10]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[10]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[10]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[10]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[11]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[11]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[11]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[11]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[11]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[11]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[11]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[12]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[12]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[12]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[12]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[12]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[12]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[12]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[13]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[13]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[13]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[13]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[13]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[13]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[13]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[14]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_address[14]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[14]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_address[14]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[14]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_address[14]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[14]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[0]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[0]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[0]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[1]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[1]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_bank[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_bank[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_bank[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_ras_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_ras_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_ras_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cas_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cas_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cas_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_we_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_we_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_we_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_cke),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_cke),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_cke),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_odt),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_odt),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_odt),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_reset_n),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_reset_n),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_reset_n),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dqs0),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(main_genericstandalone_genericstandalone_ddrphy_dqs0),
	.T(main_genericstandalone_genericstandalone_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dqs1),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(main_genericstandalone_genericstandalone_ddrphy_dqs1),
	.T(main_genericstandalone_genericstandalone_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[0]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[16]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[0]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[16]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[0]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[16]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[0]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o0),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[16]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[0]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[16]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[0]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[16]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[0]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[16]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o0),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[1]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[17]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[1]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[17]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[1]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[17]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[1]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o1),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[17]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[1]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[17]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[1]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[17]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[1]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[17]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[1])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o1),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[2]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[18]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[2]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[18]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[2]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[18]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[2]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o2),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[18]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[2]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[18]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[2]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[18]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[2]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[18]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[2])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o2),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[3]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[19]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[3]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[19]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[3]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[19]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[3]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o3),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[19]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[3]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[19]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[3]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[19]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[3]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[19]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[3])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o3),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[4]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[20]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[4]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[20]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[4]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[20]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[4]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o4),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[20]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[4]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[20]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[4]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[20]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[4]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[20]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[4])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o4),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[5]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[21]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[5]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[21]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[5]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[21]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[5]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o5),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[21]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[5]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[21]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[5]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[21]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[5]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[21]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[5])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o5),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[6]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[22]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[6]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[22]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[6]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[22]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[6]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o6),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[22]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[6]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[22]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[6]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[22]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[6]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[22]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[6])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o6),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[7]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[23]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[7]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[23]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[7]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[23]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[7]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o7),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[23]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[7]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[23]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[7]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[23]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[7]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[23]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[7])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[0] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o7),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[8]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[24]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[8]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[24]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[8]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[24]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[8]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o8),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[24]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[8]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[24]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[8]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[24]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[8]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[24]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[8])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o8),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[9]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[25]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[9]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[25]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[9]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[25]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[9]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o9),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[25]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[9]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[25]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[9]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[25]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[9]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[25]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[9])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o9),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[10]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[26]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[10]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[26]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[10]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[26]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[10]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o10),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[26]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[10]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[26]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[10]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[26]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[10]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[26]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[10])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o10),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[11]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[27]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[11]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[27]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[11]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[27]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[11]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o11),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[27]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[11]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[27]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[11]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[27]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[11]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[27]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[11])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o11),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[12]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[28]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[12]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[28]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[12]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[28]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[12]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o12),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[28]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[12]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[28]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[12]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[28]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[12]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[28]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[12])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o12),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[13]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[29]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[13]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[29]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[13]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[29]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[13]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o13),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[29]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[13]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[29]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[13]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[29]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[13]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[29]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[13])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o13),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[14]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[30]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[14]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[30]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[14]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[30]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[14]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o14),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[30]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[14]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[30]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[14]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[30]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[14]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[30]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[14])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o14),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[15]),
	.D2(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_wrdata[31]),
	.D3(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[15]),
	.D4(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_wrdata[31]),
	.D5(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[15]),
	.D6(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_wrdata[31]),
	.D7(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[15]),
	.D8(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_genericstandalone_genericstandalone_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_genericstandalone_genericstandalone_ddrphy_dq_o15),
	.TQ(main_genericstandalone_genericstandalone_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re))),
	.Q1(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[31]),
	.Q2(main_genericstandalone_genericstandalone_ddrphy_dfi_p3_rddata[15]),
	.Q3(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[31]),
	.Q4(main_genericstandalone_genericstandalone_ddrphy_dfi_p2_rddata[15]),
	.Q5(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[31]),
	.Q6(main_genericstandalone_genericstandalone_ddrphy_dfi_p1_rddata[15]),
	.Q7(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[31]),
	.Q8(main_genericstandalone_genericstandalone_ddrphy_dfi_p0_rddata[15])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((main_genericstandalone_genericstandalone_ddrphy_storage[1] & main_genericstandalone_genericstandalone_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_genericstandalone_genericstandalone_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(main_genericstandalone_genericstandalone_ddrphy_dq_o15),
	.T(main_genericstandalone_genericstandalone_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(main_genericstandalone_genericstandalone_ddrphy_dq_i_nodelay15)
);

reg [19:0] tag_mem[0:8191];
reg [12:0] memadr_1;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_tag_port_we)
		tag_mem[main_genericstandalone_genericstandalone_genericstandalone_tag_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_w;
	memadr_1 <= main_genericstandalone_genericstandalone_genericstandalone_tag_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_tag_port_dat_r = tag_mem[memadr_1];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(main_genericstandalone_genericstandalone_clk),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

assign spiflash2x_dq = main_genericstandalone_genericstandalone_spiflash_oe ? main_genericstandalone_genericstandalone_spiflash_o : 2'bz;
assign main_genericstandalone_genericstandalone_spiflash_i0 = spiflash2x_dq;

GTPE2_COMMON #(
	.PLL0_FBDIV(3'd4),
	.PLL0_FBDIV_45(3'd5),
	.PLL0_REFCLK_DIV(1'd1)
) GTPE2_COMMON (
	.BGBYPASSB(1'd1),
	.BGMONITORENB(1'd1),
	.BGPDB(1'd1),
	.BGRCALOVRD(5'd31),
	.GTREFCLK0(main_genericstandalone_genericstandalone_clk125_buf),
	.GTREFCLK1(1'd0),
	.PLL0LOCKEN(1'd1),
	.PLL0PD(1'd0),
	.PLL0REFCLKSEL(1'd1),
	.PLL0RESET(main_genericstandalone_genericstandalone_qpll_reset),
	.PLL1PD(1'd1),
	.RCALENB(1'd1),
	.PLL0LOCK(main_genericstandalone_genericstandalone_qpll_lock),
	.PLL0OUTCLK(main_genericstandalone_genericstandalone_qpll_clk),
	.PLL0OUTREFCLK(main_genericstandalone_genericstandalone_qpll_refclk)
);

GTPE2_CHANNEL #(
	.ACJTAG_DEBUG_MODE(1'd0),
	.ACJTAG_MODE(1'd0),
	.ACJTAG_RESET(1'd0),
	.ADAPT_CFG0(1'd0),
	.ALIGN_COMMA_DOUBLE("FALSE"),
	.ALIGN_COMMA_ENABLE(10'd1023),
	.ALIGN_COMMA_WORD(1'd1),
	.ALIGN_MCOMMA_DET("TRUE"),
	.ALIGN_MCOMMA_VALUE(10'd643),
	.ALIGN_PCOMMA_DET("TRUE"),
	.ALIGN_PCOMMA_VALUE(9'd380),
	.CBCC_DATA_SOURCE_SEL("ENCODED"),
	.CFOK_CFG(43'd5016522067584),
	.CFOK_CFG2(6'd32),
	.CFOK_CFG3(6'd32),
	.CFOK_CFG4(1'd0),
	.CFOK_CFG5(1'd0),
	.CFOK_CFG6(1'd0),
	.CHAN_BOND_KEEP_ALIGN("FALSE"),
	.CHAN_BOND_MAX_SKEW(1'd1),
	.CHAN_BOND_SEQ_1_1(1'd0),
	.CHAN_BOND_SEQ_1_2(1'd0),
	.CHAN_BOND_SEQ_1_3(1'd0),
	.CHAN_BOND_SEQ_1_4(1'd0),
	.CHAN_BOND_SEQ_1_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_1(1'd0),
	.CHAN_BOND_SEQ_2_2(1'd0),
	.CHAN_BOND_SEQ_2_3(1'd0),
	.CHAN_BOND_SEQ_2_4(1'd0),
	.CHAN_BOND_SEQ_2_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_USE("FALSE"),
	.CHAN_BOND_SEQ_LEN(1'd1),
	.CLK_COMMON_SWING(1'd0),
	.CLK_CORRECT_USE("FALSE"),
	.CLK_COR_KEEP_IDLE("FALSE"),
	.CLK_COR_MAX_LAT(4'd9),
	.CLK_COR_MIN_LAT(3'd7),
	.CLK_COR_PRECEDENCE("TRUE"),
	.CLK_COR_REPEAT_WAIT(1'd0),
	.CLK_COR_SEQ_1_1(9'd256),
	.CLK_COR_SEQ_1_2(1'd0),
	.CLK_COR_SEQ_1_3(1'd0),
	.CLK_COR_SEQ_1_4(1'd0),
	.CLK_COR_SEQ_1_ENABLE(4'd15),
	.CLK_COR_SEQ_2_1(9'd256),
	.CLK_COR_SEQ_2_2(1'd0),
	.CLK_COR_SEQ_2_3(1'd0),
	.CLK_COR_SEQ_2_4(1'd0),
	.CLK_COR_SEQ_2_ENABLE(4'd15),
	.CLK_COR_SEQ_2_USE("FALSE"),
	.CLK_COR_SEQ_LEN(1'd1),
	.DEC_MCOMMA_DETECT("FALSE"),
	.DEC_PCOMMA_DETECT("FALSE"),
	.DEC_VALID_COMMA_ONLY("FALSE"),
	.DMONITOR_CFG(12'd2560),
	.ES_CLK_PHASE_SEL(1'd0),
	.ES_CONTROL(1'd0),
	.ES_ERRDET_EN("FALSE"),
	.ES_EYE_SCAN_EN("FALSE"),
	.ES_HORZ_OFFSET(5'd16),
	.ES_PMA_CFG(1'd0),
	.ES_PRESCALE(1'd0),
	.ES_QUALIFIER(1'd0),
	.ES_QUAL_MASK(1'd0),
	.ES_SDATA_MASK(1'd0),
	.ES_VERT_OFFSET(1'd0),
	.FTS_DESKEW_SEQ_ENABLE(4'd15),
	.FTS_LANE_DESKEW_CFG(4'd15),
	.FTS_LANE_DESKEW_EN("FALSE"),
	.GEARBOX_MODE(1'd0),
	.LOOPBACK_CFG(1'd0),
	.OUTREFCLK_SEL_INV(2'd3),
	.PCS_PCIE_EN("FALSE"),
	.PCS_RSVD_ATTR(1'd0),
	.PD_TRANS_TIME_FROM_P2(6'd60),
	.PD_TRANS_TIME_NONE_P2(6'd60),
	.PD_TRANS_TIME_TO_P2(7'd100),
	.PMA_LOOPBACK_CFG(1'd0),
	.PMA_RSV(10'd819),
	.PMA_RSV2(14'd8256),
	.PMA_RSV3(1'd0),
	.PMA_RSV4(1'd0),
	.PMA_RSV5(1'd0),
	.PMA_RSV6(1'd0),
	.PMA_RSV7(1'd0),
	.RXBUFRESET_TIME(1'd1),
	.RXBUF_ADDR_MODE("FAST"),
	.RXBUF_EIDLE_HI_CNT(4'd8),
	.RXBUF_EIDLE_LO_CNT(1'd0),
	.RXBUF_EN("TRUE"),
	.RXBUF_RESET_ON_CB_CHANGE("TRUE"),
	.RXBUF_RESET_ON_COMMAALIGN("FALSE"),
	.RXBUF_RESET_ON_EIDLE("FALSE"),
	.RXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.RXBUF_THRESH_OVFLW(6'd61),
	.RXBUF_THRESH_OVRD("FALSE"),
	.RXBUF_THRESH_UNDFLW(3'd4),
	.RXCDRFREQRESET_TIME(1'd1),
	.RXCDRPHRESET_TIME(1'd1),
	.RXCDR_CFG(69'd314170556264376963088),
	.RXCDR_FR_RESET_ON_EIDLE(1'd0),
	.RXCDR_HOLD_DURING_EIDLE(1'd0),
	.RXCDR_LOCK_CFG(4'd9),
	.RXCDR_PH_RESET_ON_EIDLE(1'd0),
	.RXDLY_CFG(5'd31),
	.RXDLY_LCFG(6'd48),
	.RXDLY_TAP_CFG(1'd0),
	.RXGEARBOX_EN("FALSE"),
	.RXISCANRESET_TIME(1'd1),
	.RXLPMRESET_TIME(4'd15),
	.RXLPM_BIAS_STARTUP_DISABLE(1'd0),
	.RXLPM_CFG(3'd6),
	.RXLPM_CFG1(1'd0),
	.RXLPM_CM_CFG(1'd0),
	.RXLPM_GC_CFG(9'd482),
	.RXLPM_GC_CFG2(1'd1),
	.RXLPM_HF_CFG(10'd1008),
	.RXLPM_HF_CFG2(4'd10),
	.RXLPM_HF_CFG3(1'd0),
	.RXLPM_HOLD_DURING_EIDLE(1'd0),
	.RXLPM_INCM_CFG(1'd0),
	.RXLPM_IPCM_CFG(1'd1),
	.RXLPM_LF_CFG(10'd1008),
	.RXLPM_LF_CFG2(4'd10),
	.RXLPM_OSINT_CFG(3'd4),
	.RXOOB_CFG(3'd6),
	.RXOOB_CLK_CFG("PMA"),
	.RXOSCALRESET_TIME(2'd3),
	.RXOSCALRESET_TIMEOUT(1'd0),
	.RXOUT_DIV(3'd4),
	.RXPCSRESET_TIME(1'd1),
	.RXPHDLY_CFG(20'd540704),
	.RXPH_CFG(24'd12582914),
	.RXPH_MONITOR_SEL(1'd0),
	.RXPI_CFG0(1'd0),
	.RXPI_CFG1(1'd1),
	.RXPI_CFG2(1'd1),
	.RXPMARESET_TIME(2'd3),
	.RXPRBS_ERR_LOOPBACK(1'd0),
	.RXSLIDE_AUTO_WAIT(3'd7),
	.RXSLIDE_MODE("OFF"),
	.RXSYNC_MULTILANE(1'd0),
	.RXSYNC_OVRD(1'd0),
	.RXSYNC_SKIP_DA(1'd0),
	.RX_BIAS_CFG(12'd3891),
	.RX_BUFFER_CFG(1'd0),
	.RX_CLK25_DIV(3'd5),
	.RX_CLKMUX_EN(1'd1),
	.RX_CM_SEL(1'd1),
	.RX_CM_TRIM(1'd0),
	.RX_DATA_WIDTH(5'd20),
	.RX_DDI_SEL(1'd0),
	.RX_DEBUG_CFG(1'd0),
	.RX_DEFER_RESET_BUF_EN("TRUE"),
	.RX_DISPERR_SEQ_MATCH("FALSE"),
	.RX_OS_CFG(8'd128),
	.RX_SIG_VALID_DLY(4'd10),
	.RX_XCLK_SEL("RXREC"),
	.SAS_MAX_COM(7'd64),
	.SAS_MIN_COM(6'd36),
	.SATA_BURST_SEQ_LEN(3'd5),
	.SATA_BURST_VAL(3'd4),
	.SATA_EIDLE_VAL(3'd4),
	.SATA_MAX_BURST(4'd8),
	.SATA_MAX_INIT(5'd21),
	.SATA_MAX_WAKE(3'd7),
	.SATA_MIN_BURST(3'd4),
	.SATA_MIN_INIT(4'd12),
	.SATA_MIN_WAKE(3'd4),
	.SATA_PLL_CFG("VCO_3000MHZ"),
	.SHOW_REALIGN_COMMA("TRUE"),
	.SIM_RECEIVER_DETECT_PASS("TRUE"),
	.SIM_RESET_SPEEDUP("FALSE"),
	.SIM_TX_EIDLE_DRIVE_LEVEL("X"),
	.SIM_VERSION("2.0"),
	.TERM_RCAL_CFG(15'd16912),
	.TERM_RCAL_OVRD(1'd0),
	.TRANS_TIME_RATE(4'd14),
	.TST_RSV(1'd0),
	.TXBUF_EN("TRUE"),
	.TXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.TXDLY_CFG(5'd31),
	.TXDLY_LCFG(6'd48),
	.TXDLY_TAP_CFG(1'd0),
	.TXGEARBOX_EN("FALSE"),
	.TXOOB_CFG(1'd0),
	.TXOUT_DIV(3'd4),
	.TXPCSRESET_TIME(1'd1),
	.TXPHDLY_CFG(20'd540704),
	.TXPH_CFG(11'd1920),
	.TXPH_MONITOR_SEL(1'd0),
	.TXPI_CFG0(1'd0),
	.TXPI_CFG1(1'd0),
	.TXPI_CFG2(1'd0),
	.TXPI_CFG3(1'd0),
	.TXPI_CFG4(1'd0),
	.TXPI_CFG5(1'd0),
	.TXPI_GREY_SEL(1'd0),
	.TXPI_INVSTROBE_SEL(1'd0),
	.TXPI_PPMCLK_SEL("TXUSRCLK2"),
	.TXPI_PPM_CFG(1'd0),
	.TXPI_SYNFREQ_PPM(1'd1),
	.TXPMARESET_TIME(1'd1),
	.TXSYNC_MULTILANE(1'd0),
	.TXSYNC_OVRD(1'd0),
	.TXSYNC_SKIP_DA(1'd0),
	.TX_CLK25_DIV(3'd5),
	.TX_CLKMUX_EN(1'd1),
	.TX_DATA_WIDTH(5'd20),
	.TX_DEEMPH0(1'd0),
	.TX_DEEMPH1(1'd0),
	.TX_DRIVE_MODE("DIRECT"),
	.TX_EIDLE_ASSERT_DELAY(3'd6),
	.TX_EIDLE_DEASSERT_DELAY(3'd4),
	.TX_LOOPBACK_DRIVE_HIZ("FALSE"),
	.TX_MAINCURSOR_SEL(1'd0),
	.TX_MARGIN_FULL_0(7'd78),
	.TX_MARGIN_FULL_1(7'd73),
	.TX_MARGIN_FULL_2(7'd69),
	.TX_MARGIN_FULL_3(7'd66),
	.TX_MARGIN_FULL_4(7'd64),
	.TX_MARGIN_LOW_0(7'd70),
	.TX_MARGIN_LOW_1(7'd68),
	.TX_MARGIN_LOW_2(7'd66),
	.TX_MARGIN_LOW_3(7'd64),
	.TX_MARGIN_LOW_4(7'd64),
	.TX_PREDRIVER_MODE(1'd0),
	.TX_RXDETECT_CFG(13'd6194),
	.TX_RXDETECT_REF(3'd4),
	.TX_XCLK_SEL("TXOUT"),
	.UCODEER_CLR(1'd0),
	.USE_PCS_CLK_PHASE_SEL(1'd0)
) GTPE2_CHANNEL (
	.CFGRESET(1'd0),
	.CLKRSVD0(1'd0),
	.CLKRSVD1(1'd0),
	.DMONFIFORESET(1'd0),
	.DMONITORCLK(1'd0),
	.DRPADDR(main_genericstandalone_drpaddr),
	.DRPCLK(sys_clk),
	.DRPDI(main_genericstandalone_drpdi),
	.DRPEN(main_genericstandalone_drpen),
	.DRPWE(main_genericstandalone_drpwe),
	.EYESCANMODE(1'd0),
	.EYESCANRESET(1'd0),
	.EYESCANTRIGGER(1'd0),
	.GTPRXN(sfp_rxn),
	.GTPRXP(sfp_rxp),
	.GTRESETSEL(1'd0),
	.GTRSVD(1'd0),
	.GTRXRESET(main_genericstandalone_rx_reset),
	.GTTXRESET(main_genericstandalone_tx_reset),
	.LOOPBACK(1'd0),
	.PCSRSVDIN(1'd0),
	.PLL0CLK(main_genericstandalone_genericstandalone_qpll_clk),
	.PLL0REFCLK(main_genericstandalone_genericstandalone_qpll_refclk),
	.PLL1CLK(1'd0),
	.PLL1REFCLK(1'd0),
	.PMARSVDIN0(1'd0),
	.PMARSVDIN1(1'd0),
	.PMARSVDIN2(1'd0),
	.PMARSVDIN3(1'd0),
	.PMARSVDIN4(1'd0),
	.RESETOVRD(1'd0),
	.RX8B10BEN(1'd0),
	.RXADAPTSELTEST(1'd0),
	.RXBUFRESET(1'd0),
	.RXCDRFREQRESET(1'd0),
	.RXCDRHOLD(1'd0),
	.RXCDROVRDEN(1'd0),
	.RXCDRRESET(1'd0),
	.RXCDRRESETRSV(1'd0),
	.RXCHBONDEN(1'd0),
	.RXCHBONDI(1'd0),
	.RXCHBONDLEVEL(1'd0),
	.RXCHBONDMASTER(1'd0),
	.RXCHBONDSLAVE(1'd0),
	.RXCOMMADETEN(1'd0),
	.RXDDIEN(1'd0),
	.RXDFEXYDEN(1'd0),
	.RXDLYBYPASS(1'd1),
	.RXDLYEN(1'd0),
	.RXDLYOVRDEN(1'd0),
	.RXDLYSRESET(1'd0),
	.RXELECIDLEMODE(2'd3),
	.RXGEARBOXSLIP(1'd0),
	.RXLPMHFHOLD(1'd0),
	.RXLPMHFOVRDEN(1'd0),
	.RXLPMLFHOLD(1'd0),
	.RXLPMLFOVRDEN(1'd0),
	.RXLPMOSINTNTRLEN(1'd0),
	.RXLPMRESET(1'd0),
	.RXMCOMMAALIGNEN(1'd0),
	.RXOOBRESET(1'd0),
	.RXOSCALRESET(1'd0),
	.RXOSHOLD(1'd0),
	.RXOSINTCFG(2'd2),
	.RXOSINTEN(1'd1),
	.RXOSINTHOLD(1'd0),
	.RXOSINTID0(1'd0),
	.RXOSINTNTRLEN(1'd0),
	.RXOSINTOVRDEN(1'd0),
	.RXOSINTPD(1'd0),
	.RXOSINTSTROBE(1'd0),
	.RXOSINTTESTOVRDEN(1'd0),
	.RXOSOVRDEN(1'd0),
	.RXOUTCLKSEL(2'd2),
	.RXPCOMMAALIGNEN(1'd0),
	.RXPCSRESET(1'd0),
	.RXPD(1'd0),
	.RXPHALIGN(1'd0),
	.RXPHALIGNEN(1'd0),
	.RXPHDLYPD(1'd0),
	.RXPHDLYRESET(1'd0),
	.RXPHOVRDEN(1'd0),
	.RXPMARESET(1'd0),
	.RXPOLARITY(1'd0),
	.RXPRBSCNTRESET(1'd0),
	.RXPRBSSEL(1'd0),
	.RXRATE(1'd0),
	.RXRATEMODE(1'd0),
	.RXSLIDE(1'd0),
	.RXSYNCALLIN(1'd0),
	.RXSYNCIN(1'd0),
	.RXSYNCMODE(1'd0),
	.RXSYSCLKSEL(1'd0),
	.RXUSERRDY(main_genericstandalone_rx_mmcm_locked),
	.RXUSRCLK(eth_rx_half_clk),
	.RXUSRCLK2(eth_rx_half_clk),
	.SETERRSTATUS(1'd0),
	.SIGVALIDCLK(1'd0),
	.TSTIN(20'd1048575),
	.TX8B10BBYPASS(1'd0),
	.TX8B10BEN(1'd0),
	.TXBUFDIFFCTRL(3'd4),
	.TXCHARDISPMODE({main_genericstandalone_tx_data0[19], main_genericstandalone_tx_data0[9]}),
	.TXCHARDISPVAL({main_genericstandalone_tx_data0[18], main_genericstandalone_tx_data0[8]}),
	.TXCHARISK(1'd0),
	.TXCOMINIT(1'd0),
	.TXCOMSAS(1'd0),
	.TXCOMWAKE(1'd0),
	.TXDATA({main_genericstandalone_tx_data0[17:10], main_genericstandalone_tx_data0[7:0]}),
	.TXDEEMPH(1'd0),
	.TXDETECTRX(1'd0),
	.TXDIFFCTRL(4'd8),
	.TXDIFFPD(1'd0),
	.TXDLYBYPASS(1'd1),
	.TXDLYEN(1'd0),
	.TXDLYHOLD(1'd0),
	.TXDLYOVRDEN(1'd0),
	.TXDLYSRESET(1'd0),
	.TXDLYUPDOWN(1'd0),
	.TXELECIDLE(1'd0),
	.TXHEADER(1'd0),
	.TXINHIBIT(1'd0),
	.TXMAINCURSOR(1'd0),
	.TXMARGIN(1'd0),
	.TXOUTCLKSEL(2'd2),
	.TXPCSRESET(1'd0),
	.TXPD(1'd0),
	.TXPDELECIDLEMODE(1'd0),
	.TXPHALIGN(1'd0),
	.TXPHALIGNEN(1'd0),
	.TXPHDLYPD(1'd0),
	.TXPHDLYRESET(1'd0),
	.TXPHDLYTSTCLK(1'd0),
	.TXPHINIT(1'd0),
	.TXPHOVRDEN(1'd0),
	.TXPIPPMEN(1'd0),
	.TXPIPPMOVRDEN(1'd0),
	.TXPIPPMPD(1'd0),
	.TXPIPPMSEL(1'd1),
	.TXPIPPMSTEPSIZE(1'd0),
	.TXPISOPD(1'd0),
	.TXPMARESET(1'd0),
	.TXPOLARITY(1'd0),
	.TXPOSTCURSOR(1'd0),
	.TXPOSTCURSORINV(1'd0),
	.TXPRBSFORCEERR(1'd0),
	.TXPRBSSEL(1'd0),
	.TXPRECURSOR(1'd0),
	.TXPRECURSORINV(1'd0),
	.TXRATE(1'd0),
	.TXRATEMODE(1'd0),
	.TXSEQUENCE(1'd0),
	.TXSTARTSEQ(1'd0),
	.TXSWING(1'd0),
	.TXSYNCALLIN(1'd0),
	.TXSYNCIN(1'd0),
	.TXSYNCMODE(1'd0),
	.TXSYSCLKSEL(1'd0),
	.TXUSERRDY(main_genericstandalone_tx_mmcm_locked),
	.TXUSRCLK(eth_tx_half_clk),
	.TXUSRCLK2(eth_tx_half_clk),
	.DRPDO(main_genericstandalone_drpdo),
	.DRPRDY(main_genericstandalone_drprdy),
	.GTPTXN(sfp_txn),
	.GTPTXP(sfp_txp),
	.RXCHARISK({main_genericstandalone_rx_data0[18], main_genericstandalone_rx_data0[8]}),
	.RXDATA({main_genericstandalone_rx_data0[17:10], main_genericstandalone_rx_data0[7:0]}),
	.RXDISPERR({main_genericstandalone_rx_data0[19], main_genericstandalone_rx_data0[9]}),
	.RXOUTCLK(main_genericstandalone_rxoutclk),
	.RXPMARESETDONE(main_genericstandalone_rx_pma_reset_done),
	.RXRESETDONE(main_genericstandalone_rx_reset_done),
	.TXOUTCLK(main_genericstandalone_txoutclk),
	.TXRESETDONE(main_genericstandalone_tx_reset_done)
);

BUFH BUFH(
	.I(main_genericstandalone_txoutclk),
	.O(main_genericstandalone_txoutclk_rebuffer)
);

BUFG BUFG_5(
	.I(main_genericstandalone_rxoutclk),
	.O(main_genericstandalone_rxoutclk_rebuffer)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE_1 (
	.CLKFBIN(main_genericstandalone_tx_mmcm_fb),
	.CLKIN1(main_genericstandalone_txoutclk_rebuffer),
	.RST(main_genericstandalone_tx_mmcm_reset),
	.CLKFBOUT(main_genericstandalone_tx_mmcm_fb),
	.CLKOUT0(main_genericstandalone_clk_tx_half_unbuf),
	.CLKOUT1(main_genericstandalone_clk_tx_unbuf),
	.LOCKED(main_genericstandalone_tx_mmcm_locked)
);

BUFH BUFH_1(
	.I(main_genericstandalone_clk_tx_half_unbuf),
	.O(eth_tx_half_clk)
);

BUFH BUFH_2(
	.I(main_genericstandalone_clk_tx_unbuf),
	.O(eth_tx_clk)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE_2 (
	.CLKFBIN(main_genericstandalone_rx_mmcm_fb),
	.CLKIN1(main_genericstandalone_rxoutclk_rebuffer),
	.RST(main_genericstandalone_rx_mmcm_reset),
	.CLKFBOUT(main_genericstandalone_rx_mmcm_fb),
	.CLKOUT0(main_genericstandalone_clk_rx_half_unbuf),
	.CLKOUT1(main_genericstandalone_clk_rx_unbuf),
	.LOCKED(main_genericstandalone_rx_mmcm_locked)
);

BUFG BUFG_6(
	.I(main_genericstandalone_clk_rx_half_unbuf),
	.O(eth_rx_half_clk)
);

BUFG BUFG_7(
	.I(main_genericstandalone_clk_rx_unbuf),
	.O(eth_rx_clk)
);

reg [10:0] storage_2[0:4];
reg [10:0] memdat_2;
always @(posedge eth_rx_clk) begin
	if (main_genericstandalone_crc32_checker_syncfifo_wrport_we)
		storage_2[main_genericstandalone_crc32_checker_syncfifo_wrport_adr] <= main_genericstandalone_crc32_checker_syncfifo_wrport_dat_w;
	memdat_2 <= storage_2[main_genericstandalone_crc32_checker_syncfifo_wrport_adr];
end

always @(posedge eth_rx_clk) begin
end

assign main_genericstandalone_crc32_checker_syncfifo_wrport_dat_r = memdat_2;
assign main_genericstandalone_crc32_checker_syncfifo_rdport_dat_r = storage_2[main_genericstandalone_crc32_checker_syncfifo_rdport_adr];

reg [40:0] storage_3[0:63];
reg [5:0] memadr_2;
reg [5:0] memadr_3;
always @(posedge sys_clk) begin
	if (main_genericstandalone_tx_cdc_wrport_we)
		storage_3[main_genericstandalone_tx_cdc_wrport_adr] <= main_genericstandalone_tx_cdc_wrport_dat_w;
	memadr_2 <= main_genericstandalone_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memadr_3 <= main_genericstandalone_tx_cdc_rdport_adr;
end

assign main_genericstandalone_tx_cdc_wrport_dat_r = storage_3[memadr_2];
assign main_genericstandalone_tx_cdc_rdport_dat_r = storage_3[memadr_3];

reg [40:0] storage_4[0:63];
reg [5:0] memadr_4;
reg [5:0] memadr_5;
always @(posedge eth_rx_clk) begin
	if (main_genericstandalone_rx_cdc_wrport_we)
		storage_4[main_genericstandalone_rx_cdc_wrport_adr] <= main_genericstandalone_rx_cdc_wrport_dat_w;
	memadr_4 <= main_genericstandalone_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_5 <= main_genericstandalone_rx_cdc_rdport_adr;
end

assign main_genericstandalone_rx_cdc_wrport_dat_r = storage_4[memadr_4];
assign main_genericstandalone_rx_cdc_rdport_dat_r = storage_4[memadr_5];

reg [34:0] storage_5[0:3];
reg [34:0] memdat_3;
always @(posedge sys_clk) begin
	if (main_genericstandalone_writer_fifo_wrport_we)
		storage_5[main_genericstandalone_writer_fifo_wrport_adr] <= main_genericstandalone_writer_fifo_wrport_dat_w;
	memdat_3 <= storage_5[main_genericstandalone_writer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_genericstandalone_writer_fifo_wrport_dat_r = memdat_3;
assign main_genericstandalone_writer_fifo_rdport_dat_r = storage_5[main_genericstandalone_writer_fifo_rdport_adr];

reg [31:0] mem_1[0:381];
reg [8:0] memadr_6;
reg [8:0] memadr_7;
always @(posedge sys_clk) begin
	if (main_genericstandalone_writer_memory0_we)
		mem_1[main_genericstandalone_writer_memory0_adr] <= main_genericstandalone_writer_memory0_dat_w;
	memadr_6 <= main_genericstandalone_writer_memory0_adr;
end

always @(posedge sys_clk) begin
	memadr_7 <= main_genericstandalone_sram0_adr0;
end

assign main_genericstandalone_writer_memory0_dat_r = mem_1[memadr_6];
assign main_genericstandalone_sram0_dat_r0 = mem_1[memadr_7];

reg [31:0] mem_2[0:381];
reg [8:0] memadr_8;
reg [8:0] memadr_9;
always @(posedge sys_clk) begin
	if (main_genericstandalone_writer_memory1_we)
		mem_2[main_genericstandalone_writer_memory1_adr] <= main_genericstandalone_writer_memory1_dat_w;
	memadr_8 <= main_genericstandalone_writer_memory1_adr;
end

always @(posedge sys_clk) begin
	memadr_9 <= main_genericstandalone_sram1_adr0;
end

assign main_genericstandalone_writer_memory1_dat_r = mem_2[memadr_8];
assign main_genericstandalone_sram1_dat_r0 = mem_2[memadr_9];

reg [31:0] mem_3[0:381];
reg [8:0] memadr_10;
reg [8:0] memadr_11;
always @(posedge sys_clk) begin
	if (main_genericstandalone_writer_memory2_we)
		mem_3[main_genericstandalone_writer_memory2_adr] <= main_genericstandalone_writer_memory2_dat_w;
	memadr_10 <= main_genericstandalone_writer_memory2_adr;
end

always @(posedge sys_clk) begin
	memadr_11 <= main_genericstandalone_sram2_adr0;
end

assign main_genericstandalone_writer_memory2_dat_r = mem_3[memadr_10];
assign main_genericstandalone_sram2_dat_r0 = mem_3[memadr_11];

reg [31:0] mem_4[0:381];
reg [8:0] memadr_12;
reg [8:0] memadr_13;
always @(posedge sys_clk) begin
	if (main_genericstandalone_writer_memory3_we)
		mem_4[main_genericstandalone_writer_memory3_adr] <= main_genericstandalone_writer_memory3_dat_w;
	memadr_12 <= main_genericstandalone_writer_memory3_adr;
end

always @(posedge sys_clk) begin
	memadr_13 <= main_genericstandalone_sram3_adr0;
end

assign main_genericstandalone_writer_memory3_dat_r = mem_4[memadr_12];
assign main_genericstandalone_sram3_dat_r0 = mem_4[memadr_13];

reg [13:0] storage_6[0:3];
reg [13:0] memdat_4;
always @(posedge sys_clk) begin
	if (main_genericstandalone_reader_fifo_wrport_we)
		storage_6[main_genericstandalone_reader_fifo_wrport_adr] <= main_genericstandalone_reader_fifo_wrport_dat_w;
	memdat_4 <= storage_6[main_genericstandalone_reader_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_genericstandalone_reader_fifo_wrport_dat_r = memdat_4;
assign main_genericstandalone_reader_fifo_rdport_dat_r = storage_6[main_genericstandalone_reader_fifo_rdport_adr];

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(31'd1082130432)
) mor1kx_1 (
	.clk(sys_kernel_clk),
	.dwbm_ack_i(main_genericstandalone_kernel_cpu_dbus_ack),
	.dwbm_dat_i(main_genericstandalone_kernel_cpu_dbus_dat_r),
	.dwbm_err_i(main_genericstandalone_kernel_cpu_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(main_genericstandalone_kernel_cpu_interrupt),
	.iwbm_ack_i(main_genericstandalone_kernel_cpu_ibus_ack),
	.iwbm_dat_i(main_genericstandalone_kernel_cpu_ibus_dat_r),
	.iwbm_err_i(main_genericstandalone_kernel_cpu_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_kernel_rst),
	.dwbm_adr_o(main_genericstandalone_kernel_cpu_d_adr_o),
	.dwbm_bte_o(main_genericstandalone_kernel_cpu_dbus_bte),
	.dwbm_cti_o(main_genericstandalone_kernel_cpu_dbus_cti),
	.dwbm_cyc_o(main_genericstandalone_kernel_cpu_dbus_cyc),
	.dwbm_dat_o(main_genericstandalone_kernel_cpu_dbus_dat_w),
	.dwbm_sel_o(main_genericstandalone_kernel_cpu_dbus_sel),
	.dwbm_stb_o(main_genericstandalone_kernel_cpu_dbus_stb),
	.dwbm_we_o(main_genericstandalone_kernel_cpu_dbus_we),
	.iwbm_adr_o(main_genericstandalone_kernel_cpu_i_adr_o),
	.iwbm_bte_o(main_genericstandalone_kernel_cpu_ibus_bte),
	.iwbm_cti_o(main_genericstandalone_kernel_cpu_ibus_cti),
	.iwbm_cyc_o(main_genericstandalone_kernel_cpu_ibus_cyc),
	.iwbm_dat_o(main_genericstandalone_kernel_cpu_ibus_dat_w),
	.iwbm_sel_o(main_genericstandalone_kernel_cpu_ibus_sel),
	.iwbm_stb_o(main_genericstandalone_kernel_cpu_ibus_stb),
	.iwbm_we_o(main_genericstandalone_kernel_cpu_ibus_we)
);

reg [7:0] mem_5[0:37];
reg [5:0] memadr_14;
always @(posedge sys_clk) begin
	memadr_14 <= main_add_identifier_adr;
end

assign main_add_identifier_dat_r = mem_5[memadr_14];

initial begin
	$readmemh("mem_5.init", mem_5);
end

assign i2c_scl = main_i2c_tstriple0_oe ? main_i2c_tstriple0_o : 1'bz;
assign main_i2c_tstriple0_i = i2c_scl;

assign i2c_sda = main_i2c_tstriple1_oe ? main_i2c_tstriple1_o : 1'bz;
assign main_i2c_tstriple1_i = i2c_sda;

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_16 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x0_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x0_serdes_i1[7]),
	.Q2(main_inout_8x0_serdes_i1[6]),
	.Q3(main_inout_8x0_serdes_i1[5]),
	.Q4(main_inout_8x0_serdes_i1[4]),
	.Q5(main_inout_8x0_serdes_i1[3]),
	.Q6(main_inout_8x0_serdes_i1[2]),
	.Q7(main_inout_8x0_serdes_i1[1]),
	.Q8(main_inout_8x0_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x0_serdes_o1[0]),
	.D2(main_inout_8x0_serdes_o1[1]),
	.D3(main_inout_8x0_serdes_o1[2]),
	.D4(main_inout_8x0_serdes_o1[3]),
	.D5(main_inout_8x0_serdes_o1[4]),
	.D6(main_inout_8x0_serdes_o1[5]),
	.D7(main_inout_8x0_serdes_o1[6]),
	.D8(main_inout_8x0_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x0_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x0_serdes_pad_o1),
	.TQ(main_inout_8x0_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE (
	.I(main_inout_8x0_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x0_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x0_serdes_t_out)),
	.T(main_inout_8x0_serdes_t_out),
	.IO(dio0_p),
	.IOB(dio0_n),
	.O(main_inout_8x0_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_17 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x1_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x1_serdes_i1[7]),
	.Q2(main_inout_8x1_serdes_i1[6]),
	.Q3(main_inout_8x1_serdes_i1[5]),
	.Q4(main_inout_8x1_serdes_i1[4]),
	.Q5(main_inout_8x1_serdes_i1[3]),
	.Q6(main_inout_8x1_serdes_i1[2]),
	.Q7(main_inout_8x1_serdes_i1[1]),
	.Q8(main_inout_8x1_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x1_serdes_o1[0]),
	.D2(main_inout_8x1_serdes_o1[1]),
	.D3(main_inout_8x1_serdes_o1[2]),
	.D4(main_inout_8x1_serdes_o1[3]),
	.D5(main_inout_8x1_serdes_o1[4]),
	.D6(main_inout_8x1_serdes_o1[5]),
	.D7(main_inout_8x1_serdes_o1[6]),
	.D8(main_inout_8x1_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x1_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x1_serdes_pad_o1),
	.TQ(main_inout_8x1_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_1 (
	.I(main_inout_8x1_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x1_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x1_serdes_t_out)),
	.T(main_inout_8x1_serdes_t_out),
	.IO(dio0_p_1),
	.IOB(dio0_n_1),
	.O(main_inout_8x1_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_18 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x2_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x2_serdes_i1[7]),
	.Q2(main_inout_8x2_serdes_i1[6]),
	.Q3(main_inout_8x2_serdes_i1[5]),
	.Q4(main_inout_8x2_serdes_i1[4]),
	.Q5(main_inout_8x2_serdes_i1[3]),
	.Q6(main_inout_8x2_serdes_i1[2]),
	.Q7(main_inout_8x2_serdes_i1[1]),
	.Q8(main_inout_8x2_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x2_serdes_o1[0]),
	.D2(main_inout_8x2_serdes_o1[1]),
	.D3(main_inout_8x2_serdes_o1[2]),
	.D4(main_inout_8x2_serdes_o1[3]),
	.D5(main_inout_8x2_serdes_o1[4]),
	.D6(main_inout_8x2_serdes_o1[5]),
	.D7(main_inout_8x2_serdes_o1[6]),
	.D8(main_inout_8x2_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x2_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x2_serdes_pad_o1),
	.TQ(main_inout_8x2_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_2 (
	.I(main_inout_8x2_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x2_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x2_serdes_t_out)),
	.T(main_inout_8x2_serdes_t_out),
	.IO(dio0_p_2),
	.IOB(dio0_n_2),
	.O(main_inout_8x2_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_19 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x3_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x3_serdes_i1[7]),
	.Q2(main_inout_8x3_serdes_i1[6]),
	.Q3(main_inout_8x3_serdes_i1[5]),
	.Q4(main_inout_8x3_serdes_i1[4]),
	.Q5(main_inout_8x3_serdes_i1[3]),
	.Q6(main_inout_8x3_serdes_i1[2]),
	.Q7(main_inout_8x3_serdes_i1[1]),
	.Q8(main_inout_8x3_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x3_serdes_o1[0]),
	.D2(main_inout_8x3_serdes_o1[1]),
	.D3(main_inout_8x3_serdes_o1[2]),
	.D4(main_inout_8x3_serdes_o1[3]),
	.D5(main_inout_8x3_serdes_o1[4]),
	.D6(main_inout_8x3_serdes_o1[5]),
	.D7(main_inout_8x3_serdes_o1[6]),
	.D8(main_inout_8x3_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x3_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x3_serdes_pad_o1),
	.TQ(main_inout_8x3_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_3 (
	.I(main_inout_8x3_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x3_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x3_serdes_t_out)),
	.T(main_inout_8x3_serdes_t_out),
	.IO(dio0_p_3),
	.IOB(dio0_n_3),
	.O(main_inout_8x3_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_20 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x4_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x4_serdes_i1[7]),
	.Q2(main_inout_8x4_serdes_i1[6]),
	.Q3(main_inout_8x4_serdes_i1[5]),
	.Q4(main_inout_8x4_serdes_i1[4]),
	.Q5(main_inout_8x4_serdes_i1[3]),
	.Q6(main_inout_8x4_serdes_i1[2]),
	.Q7(main_inout_8x4_serdes_i1[1]),
	.Q8(main_inout_8x4_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x4_serdes_o1[0]),
	.D2(main_inout_8x4_serdes_o1[1]),
	.D3(main_inout_8x4_serdes_o1[2]),
	.D4(main_inout_8x4_serdes_o1[3]),
	.D5(main_inout_8x4_serdes_o1[4]),
	.D6(main_inout_8x4_serdes_o1[5]),
	.D7(main_inout_8x4_serdes_o1[6]),
	.D8(main_inout_8x4_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x4_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x4_serdes_pad_o1),
	.TQ(main_inout_8x4_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_4 (
	.I(main_inout_8x4_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x4_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x4_serdes_t_out)),
	.T(main_inout_8x4_serdes_t_out),
	.IO(dio0_p_4),
	.IOB(dio0_n_4),
	.O(main_inout_8x4_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_21 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x5_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x5_serdes_i1[7]),
	.Q2(main_inout_8x5_serdes_i1[6]),
	.Q3(main_inout_8x5_serdes_i1[5]),
	.Q4(main_inout_8x5_serdes_i1[4]),
	.Q5(main_inout_8x5_serdes_i1[3]),
	.Q6(main_inout_8x5_serdes_i1[2]),
	.Q7(main_inout_8x5_serdes_i1[1]),
	.Q8(main_inout_8x5_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x5_serdes_o1[0]),
	.D2(main_inout_8x5_serdes_o1[1]),
	.D3(main_inout_8x5_serdes_o1[2]),
	.D4(main_inout_8x5_serdes_o1[3]),
	.D5(main_inout_8x5_serdes_o1[4]),
	.D6(main_inout_8x5_serdes_o1[5]),
	.D7(main_inout_8x5_serdes_o1[6]),
	.D8(main_inout_8x5_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x5_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x5_serdes_pad_o1),
	.TQ(main_inout_8x5_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_5 (
	.I(main_inout_8x5_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x5_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x5_serdes_t_out)),
	.T(main_inout_8x5_serdes_t_out),
	.IO(dio0_p_5),
	.IOB(dio0_n_5),
	.O(main_inout_8x5_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_22 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x6_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x6_serdes_i1[7]),
	.Q2(main_inout_8x6_serdes_i1[6]),
	.Q3(main_inout_8x6_serdes_i1[5]),
	.Q4(main_inout_8x6_serdes_i1[4]),
	.Q5(main_inout_8x6_serdes_i1[3]),
	.Q6(main_inout_8x6_serdes_i1[2]),
	.Q7(main_inout_8x6_serdes_i1[1]),
	.Q8(main_inout_8x6_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x6_serdes_o1[0]),
	.D2(main_inout_8x6_serdes_o1[1]),
	.D3(main_inout_8x6_serdes_o1[2]),
	.D4(main_inout_8x6_serdes_o1[3]),
	.D5(main_inout_8x6_serdes_o1[4]),
	.D6(main_inout_8x6_serdes_o1[5]),
	.D7(main_inout_8x6_serdes_o1[6]),
	.D8(main_inout_8x6_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x6_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x6_serdes_pad_o1),
	.TQ(main_inout_8x6_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_6 (
	.I(main_inout_8x6_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x6_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x6_serdes_t_out)),
	.T(main_inout_8x6_serdes_t_out),
	.IO(dio0_p_6),
	.IOB(dio0_n_6),
	.O(main_inout_8x6_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_23 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x7_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x7_serdes_i1[7]),
	.Q2(main_inout_8x7_serdes_i1[6]),
	.Q3(main_inout_8x7_serdes_i1[5]),
	.Q4(main_inout_8x7_serdes_i1[4]),
	.Q5(main_inout_8x7_serdes_i1[3]),
	.Q6(main_inout_8x7_serdes_i1[2]),
	.Q7(main_inout_8x7_serdes_i1[1]),
	.Q8(main_inout_8x7_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_inout_8x7_serdes_o1[0]),
	.D2(main_inout_8x7_serdes_o1[1]),
	.D3(main_inout_8x7_serdes_o1[2]),
	.D4(main_inout_8x7_serdes_o1[3]),
	.D5(main_inout_8x7_serdes_o1[4]),
	.D6(main_inout_8x7_serdes_o1[5]),
	.D7(main_inout_8x7_serdes_o1[6]),
	.D8(main_inout_8x7_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x7_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x7_serdes_pad_o1),
	.TQ(main_inout_8x7_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_7 (
	.I(main_inout_8x7_serdes_pad_o0),
	.IBUFDISABLE((~main_inout_8x7_serdes_t_out)),
	.INTERMDISABLE((~main_inout_8x7_serdes_t_out)),
	.T(main_inout_8x7_serdes_t_out),
	.IO(dio0_p_7),
	.IOB(dio0_n_7),
	.O(main_inout_8x7_serdes_pad_i0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_53 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x0_o[0]),
	.D2(main_output_8x0_o[1]),
	.D3(main_output_8x0_o[2]),
	.D4(main_output_8x0_o[3]),
	.D5(main_output_8x0_o[4]),
	.D6(main_output_8x0_o[5]),
	.D7(main_output_8x0_o[6]),
	.D8(main_output_8x0_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x0_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x0_pad_o),
	.TQ(main_output_8x0_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_8 (
	.I(main_output_8x0_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x0_t_out),
	.IO(dio1_p),
	.IOB(dio1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_54 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x1_o[0]),
	.D2(main_output_8x1_o[1]),
	.D3(main_output_8x1_o[2]),
	.D4(main_output_8x1_o[3]),
	.D5(main_output_8x1_o[4]),
	.D6(main_output_8x1_o[5]),
	.D7(main_output_8x1_o[6]),
	.D8(main_output_8x1_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x1_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x1_pad_o),
	.TQ(main_output_8x1_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_9 (
	.I(main_output_8x1_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x1_t_out),
	.IO(dio1_p_1),
	.IOB(dio1_n_1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_55 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x2_o[0]),
	.D2(main_output_8x2_o[1]),
	.D3(main_output_8x2_o[2]),
	.D4(main_output_8x2_o[3]),
	.D5(main_output_8x2_o[4]),
	.D6(main_output_8x2_o[5]),
	.D7(main_output_8x2_o[6]),
	.D8(main_output_8x2_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x2_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x2_pad_o),
	.TQ(main_output_8x2_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_10 (
	.I(main_output_8x2_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x2_t_out),
	.IO(dio1_p_2),
	.IOB(dio1_n_2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_56 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x3_o[0]),
	.D2(main_output_8x3_o[1]),
	.D3(main_output_8x3_o[2]),
	.D4(main_output_8x3_o[3]),
	.D5(main_output_8x3_o[4]),
	.D6(main_output_8x3_o[5]),
	.D7(main_output_8x3_o[6]),
	.D8(main_output_8x3_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x3_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x3_pad_o),
	.TQ(main_output_8x3_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_11 (
	.I(main_output_8x3_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x3_t_out),
	.IO(dio1_p_3),
	.IOB(dio1_n_3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_57 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x4_o[0]),
	.D2(main_output_8x4_o[1]),
	.D3(main_output_8x4_o[2]),
	.D4(main_output_8x4_o[3]),
	.D5(main_output_8x4_o[4]),
	.D6(main_output_8x4_o[5]),
	.D7(main_output_8x4_o[6]),
	.D8(main_output_8x4_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x4_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x4_pad_o),
	.TQ(main_output_8x4_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_12 (
	.I(main_output_8x4_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x4_t_out),
	.IO(dio1_p_4),
	.IOB(dio1_n_4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_58 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x5_o[0]),
	.D2(main_output_8x5_o[1]),
	.D3(main_output_8x5_o[2]),
	.D4(main_output_8x5_o[3]),
	.D5(main_output_8x5_o[4]),
	.D6(main_output_8x5_o[5]),
	.D7(main_output_8x5_o[6]),
	.D8(main_output_8x5_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x5_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x5_pad_o),
	.TQ(main_output_8x5_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_13 (
	.I(main_output_8x5_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x5_t_out),
	.IO(dio1_p_5),
	.IOB(dio1_n_5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_59 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x6_o[0]),
	.D2(main_output_8x6_o[1]),
	.D3(main_output_8x6_o[2]),
	.D4(main_output_8x6_o[3]),
	.D5(main_output_8x6_o[4]),
	.D6(main_output_8x6_o[5]),
	.D7(main_output_8x6_o[6]),
	.D8(main_output_8x6_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x6_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x6_pad_o),
	.TQ(main_output_8x6_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_14 (
	.I(main_output_8x6_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x6_t_out),
	.IO(dio1_p_6),
	.IOB(dio1_n_6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_60 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x7_o[0]),
	.D2(main_output_8x7_o[1]),
	.D3(main_output_8x7_o[2]),
	.D4(main_output_8x7_o[3]),
	.D5(main_output_8x7_o[4]),
	.D6(main_output_8x7_o[5]),
	.D7(main_output_8x7_o[6]),
	.D8(main_output_8x7_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x7_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x7_pad_o),
	.TQ(main_output_8x7_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_15 (
	.I(main_output_8x7_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x7_t_out),
	.IO(dio1_p_7),
	.IOB(dio1_n_7)
);

OBUFTDS OBUFTDS_2(
	.I(main_spimaster0_interface_cs1[0]),
	.T(main_spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[0]),
	.OB(urukul2_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_3(
	.I(main_spimaster0_interface_cs1[1]),
	.T(main_spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[1]),
	.OB(urukul2_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_4(
	.I(main_spimaster0_interface_cs1[2]),
	.T(main_spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[2]),
	.OB(urukul2_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_5(
	.I(main_spimaster0_interface_clk),
	.T(main_spimaster0_interface_offline),
	.O(urukul2_spi_p_clk),
	.OB(urukul2_spi_n_clk)
);

IOBUFDS IOBUFDS(
	.I(main_spimaster0_interface_sdo),
	.T((main_spimaster0_interface_offline | main_spimaster0_interface_half_duplex)),
	.IO(urukul2_spi_p_mosi),
	.IOB(urukul2_spi_n_mosi),
	.O(main_spimaster0_interface_mosi)
);

IOBUFDS IOBUFDS_1(
	.I(main_spimaster0_interface_sdo),
	.T(1'd1),
	.IO(urukul2_spi_p_miso),
	.IOB(urukul2_spi_n_miso),
	.O(main_spimaster0_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_61 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x8_o[0]),
	.D2(main_output_8x8_o[1]),
	.D3(main_output_8x8_o[2]),
	.D4(main_output_8x8_o[3]),
	.D5(main_output_8x8_o[4]),
	.D6(main_output_8x8_o[5]),
	.D7(main_output_8x8_o[6]),
	.D8(main_output_8x8_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x8_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x8_pad_o),
	.TQ(main_output_8x8_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_16 (
	.I(main_output_8x8_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x8_t_out),
	.IO(urukul2_io_update_p),
	.IOB(urukul2_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_62 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x9_o[0]),
	.D2(main_output_8x9_o[1]),
	.D3(main_output_8x9_o[2]),
	.D4(main_output_8x9_o[3]),
	.D5(main_output_8x9_o[4]),
	.D6(main_output_8x9_o[5]),
	.D7(main_output_8x9_o[6]),
	.D8(main_output_8x9_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x9_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x9_pad_o),
	.TQ(main_output_8x9_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_17 (
	.I(main_output_8x9_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x9_t_out),
	.IO(urukul2_sw0_p),
	.IOB(urukul2_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_63 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x10_o[0]),
	.D2(main_output_8x10_o[1]),
	.D3(main_output_8x10_o[2]),
	.D4(main_output_8x10_o[3]),
	.D5(main_output_8x10_o[4]),
	.D6(main_output_8x10_o[5]),
	.D7(main_output_8x10_o[6]),
	.D8(main_output_8x10_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x10_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x10_pad_o),
	.TQ(main_output_8x10_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_18 (
	.I(main_output_8x10_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x10_t_out),
	.IO(urukul2_sw1_p),
	.IOB(urukul2_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_64 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x11_o[0]),
	.D2(main_output_8x11_o[1]),
	.D3(main_output_8x11_o[2]),
	.D4(main_output_8x11_o[3]),
	.D5(main_output_8x11_o[4]),
	.D6(main_output_8x11_o[5]),
	.D7(main_output_8x11_o[6]),
	.D8(main_output_8x11_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x11_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x11_pad_o),
	.TQ(main_output_8x11_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_19 (
	.I(main_output_8x11_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x11_t_out),
	.IO(urukul2_sw2_p),
	.IOB(urukul2_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_65 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x12_o[0]),
	.D2(main_output_8x12_o[1]),
	.D3(main_output_8x12_o[2]),
	.D4(main_output_8x12_o[3]),
	.D5(main_output_8x12_o[4]),
	.D6(main_output_8x12_o[5]),
	.D7(main_output_8x12_o[6]),
	.D8(main_output_8x12_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x12_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x12_pad_o),
	.TQ(main_output_8x12_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_20 (
	.I(main_output_8x12_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x12_t_out),
	.IO(urukul2_sw3_p),
	.IOB(urukul2_sw3_n)
);

OBUFTDS OBUFTDS_6(
	.I(main_spimaster1_interface_cs1[0]),
	.T(main_spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[0]),
	.OB(urukul4_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_7(
	.I(main_spimaster1_interface_cs1[1]),
	.T(main_spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[1]),
	.OB(urukul4_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_8(
	.I(main_spimaster1_interface_cs1[2]),
	.T(main_spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[2]),
	.OB(urukul4_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_9(
	.I(main_spimaster1_interface_clk),
	.T(main_spimaster1_interface_offline),
	.O(urukul4_spi_p_clk),
	.OB(urukul4_spi_n_clk)
);

IOBUFDS IOBUFDS_2(
	.I(main_spimaster1_interface_sdo),
	.T((main_spimaster1_interface_offline | main_spimaster1_interface_half_duplex)),
	.IO(urukul4_spi_p_mosi),
	.IOB(urukul4_spi_n_mosi),
	.O(main_spimaster1_interface_mosi)
);

IOBUFDS IOBUFDS_3(
	.I(main_spimaster1_interface_sdo),
	.T(1'd1),
	.IO(urukul4_spi_p_miso),
	.IOB(urukul4_spi_n_miso),
	.O(main_spimaster1_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_66 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x13_o[0]),
	.D2(main_output_8x13_o[1]),
	.D3(main_output_8x13_o[2]),
	.D4(main_output_8x13_o[3]),
	.D5(main_output_8x13_o[4]),
	.D6(main_output_8x13_o[5]),
	.D7(main_output_8x13_o[6]),
	.D8(main_output_8x13_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x13_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x13_pad_o),
	.TQ(main_output_8x13_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_21 (
	.I(main_output_8x13_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x13_t_out),
	.IO(urukul4_io_update_p),
	.IOB(urukul4_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_67 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x14_o[0]),
	.D2(main_output_8x14_o[1]),
	.D3(main_output_8x14_o[2]),
	.D4(main_output_8x14_o[3]),
	.D5(main_output_8x14_o[4]),
	.D6(main_output_8x14_o[5]),
	.D7(main_output_8x14_o[6]),
	.D8(main_output_8x14_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x14_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x14_pad_o),
	.TQ(main_output_8x14_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_22 (
	.I(main_output_8x14_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x14_t_out),
	.IO(urukul4_sw0_p),
	.IOB(urukul4_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_68 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x15_o[0]),
	.D2(main_output_8x15_o[1]),
	.D3(main_output_8x15_o[2]),
	.D4(main_output_8x15_o[3]),
	.D5(main_output_8x15_o[4]),
	.D6(main_output_8x15_o[5]),
	.D7(main_output_8x15_o[6]),
	.D8(main_output_8x15_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x15_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x15_pad_o),
	.TQ(main_output_8x15_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_23 (
	.I(main_output_8x15_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x15_t_out),
	.IO(urukul4_sw1_p),
	.IOB(urukul4_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_69 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x16_o[0]),
	.D2(main_output_8x16_o[1]),
	.D3(main_output_8x16_o[2]),
	.D4(main_output_8x16_o[3]),
	.D5(main_output_8x16_o[4]),
	.D6(main_output_8x16_o[5]),
	.D7(main_output_8x16_o[6]),
	.D8(main_output_8x16_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x16_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x16_pad_o),
	.TQ(main_output_8x16_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_24 (
	.I(main_output_8x16_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x16_t_out),
	.IO(urukul4_sw2_p),
	.IOB(urukul4_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_70 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x17_o[0]),
	.D2(main_output_8x17_o[1]),
	.D3(main_output_8x17_o[2]),
	.D4(main_output_8x17_o[3]),
	.D5(main_output_8x17_o[4]),
	.D6(main_output_8x17_o[5]),
	.D7(main_output_8x17_o[6]),
	.D8(main_output_8x17_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x17_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x17_pad_o),
	.TQ(main_output_8x17_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_25 (
	.I(main_output_8x17_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x17_t_out),
	.IO(urukul4_sw3_p),
	.IOB(urukul4_sw3_n)
);

OBUFTDS OBUFTDS_10(
	.I(main_spimaster2_interface_cs1[0]),
	.T(main_spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[0]),
	.OB(urukul6_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_11(
	.I(main_spimaster2_interface_cs1[1]),
	.T(main_spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[1]),
	.OB(urukul6_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_12(
	.I(main_spimaster2_interface_cs1[2]),
	.T(main_spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[2]),
	.OB(urukul6_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_13(
	.I(main_spimaster2_interface_clk),
	.T(main_spimaster2_interface_offline),
	.O(urukul6_spi_p_clk),
	.OB(urukul6_spi_n_clk)
);

IOBUFDS IOBUFDS_4(
	.I(main_spimaster2_interface_sdo),
	.T((main_spimaster2_interface_offline | main_spimaster2_interface_half_duplex)),
	.IO(urukul6_spi_p_mosi),
	.IOB(urukul6_spi_n_mosi),
	.O(main_spimaster2_interface_mosi)
);

IOBUFDS IOBUFDS_5(
	.I(main_spimaster2_interface_sdo),
	.T(1'd1),
	.IO(urukul6_spi_p_miso),
	.IOB(urukul6_spi_n_miso),
	.O(main_spimaster2_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_71 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x18_o[0]),
	.D2(main_output_8x18_o[1]),
	.D3(main_output_8x18_o[2]),
	.D4(main_output_8x18_o[3]),
	.D5(main_output_8x18_o[4]),
	.D6(main_output_8x18_o[5]),
	.D7(main_output_8x18_o[6]),
	.D8(main_output_8x18_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x18_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x18_pad_o),
	.TQ(main_output_8x18_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_26 (
	.I(main_output_8x18_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x18_t_out),
	.IO(urukul6_io_update_p),
	.IOB(urukul6_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_72 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x19_o[0]),
	.D2(main_output_8x19_o[1]),
	.D3(main_output_8x19_o[2]),
	.D4(main_output_8x19_o[3]),
	.D5(main_output_8x19_o[4]),
	.D6(main_output_8x19_o[5]),
	.D7(main_output_8x19_o[6]),
	.D8(main_output_8x19_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x19_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x19_pad_o),
	.TQ(main_output_8x19_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_27 (
	.I(main_output_8x19_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x19_t_out),
	.IO(urukul6_sw0_p),
	.IOB(urukul6_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_73 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x20_o[0]),
	.D2(main_output_8x20_o[1]),
	.D3(main_output_8x20_o[2]),
	.D4(main_output_8x20_o[3]),
	.D5(main_output_8x20_o[4]),
	.D6(main_output_8x20_o[5]),
	.D7(main_output_8x20_o[6]),
	.D8(main_output_8x20_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x20_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x20_pad_o),
	.TQ(main_output_8x20_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_28 (
	.I(main_output_8x20_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x20_t_out),
	.IO(urukul6_sw1_p),
	.IOB(urukul6_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_74 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x21_o[0]),
	.D2(main_output_8x21_o[1]),
	.D3(main_output_8x21_o[2]),
	.D4(main_output_8x21_o[3]),
	.D5(main_output_8x21_o[4]),
	.D6(main_output_8x21_o[5]),
	.D7(main_output_8x21_o[6]),
	.D8(main_output_8x21_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x21_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x21_pad_o),
	.TQ(main_output_8x21_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_29 (
	.I(main_output_8x21_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x21_t_out),
	.IO(urukul6_sw2_p),
	.IOB(urukul6_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_75 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(main_output_8x22_o[0]),
	.D2(main_output_8x22_o[1]),
	.D3(main_output_8x22_o[2]),
	.D4(main_output_8x22_o[3]),
	.D5(main_output_8x22_o[4]),
	.D6(main_output_8x22_o[5]),
	.D7(main_output_8x22_o[6]),
	.D8(main_output_8x22_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x22_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x22_pad_o),
	.TQ(main_output_8x22_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_30 (
	.I(main_output_8x22_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(main_output_8x22_t_out),
	.IO(urukul6_sw3_p),
	.IOB(urukul6_sw3_n)
);

IBUFGDS #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("FALSE")
) IBUFGDS (
	.I(si5324_clkout_fabric_p),
	.IB(si5324_clkout_fabric_n),
	.O(main_rtio_crg_clk_synth_se)
);

PLLE2_ADV #(
	.BANDWIDTH("HIGH"),
	.CLKFBOUT_MULT(4'd12),
	.CLKIN1_PERIOD(8.0),
	.CLKIN2_PERIOD(8.0),
	.CLKOUT0_DIVIDE(2'd3),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd12),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.001),
	.STARTUP_WAIT("FALSE")
) PLLE2_ADV (
	.CLKFBIN(main_rtio_crg_fb_clk),
	.CLKIN2(main_rtio_crg_clk_synth_se),
	.CLKINSEL(1'd0),
	.RST(main_rtio_crg_storage),
	.CLKFBOUT(main_rtio_crg_fb_clk),
	.CLKOUT0(main_rtio_crg_rtiox4_clk),
	.CLKOUT1(main_rtio_crg_rtio_clk),
	.LOCKED(main_rtio_crg_pll_locked)
);

BUFG BUFG_8(
	.I(main_rtio_crg_rtio_clk),
	.O(rtio_clk)
);

BUFG BUFG_9(
	.I(main_rtio_crg_rtiox4_clk),
	.O(rtiox4_clk)
);

reg [13:0] latency_compensation[0:36];
reg [5:0] memadr_15;
always @(posedge rsys_clk) begin
	memadr_15 <= main_rtio_core_outputs_lanedistributor_adr;
end

assign main_rtio_core_outputs_lanedistributor_dat_r = latency_compensation[memadr_15];

initial begin
	$readmemh("latency_compensation.init", latency_compensation);
end

reg [115:0] storage_7[0:127];
reg [6:0] memadr_16;
reg [6:0] memadr_17;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered0_wrport_we)
		storage_7[main_rtio_core_outputs_asyncfifobuffered0_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
	memadr_16 <= main_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_17 <= main_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r = storage_7[memadr_16];
assign main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r = storage_7[memadr_17];

reg [115:0] storage_8[0:127];
reg [6:0] memadr_18;
reg [6:0] memadr_19;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered1_wrport_we)
		storage_8[main_rtio_core_outputs_asyncfifobuffered1_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
	memadr_18 <= main_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_19 <= main_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r = storage_8[memadr_18];
assign main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r = storage_8[memadr_19];

reg [115:0] storage_9[0:127];
reg [6:0] memadr_20;
reg [6:0] memadr_21;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered2_wrport_we)
		storage_9[main_rtio_core_outputs_asyncfifobuffered2_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
	memadr_20 <= main_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_21 <= main_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r = storage_9[memadr_20];
assign main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r = storage_9[memadr_21];

reg [115:0] storage_10[0:127];
reg [6:0] memadr_22;
reg [6:0] memadr_23;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered3_wrport_we)
		storage_10[main_rtio_core_outputs_asyncfifobuffered3_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
	memadr_22 <= main_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_23 <= main_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r = storage_10[memadr_22];
assign main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r = storage_10[memadr_23];

reg [115:0] storage_11[0:127];
reg [6:0] memadr_24;
reg [6:0] memadr_25;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered4_wrport_we)
		storage_11[main_rtio_core_outputs_asyncfifobuffered4_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
	memadr_24 <= main_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_25 <= main_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r = storage_11[memadr_24];
assign main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r = storage_11[memadr_25];

reg [115:0] storage_12[0:127];
reg [6:0] memadr_26;
reg [6:0] memadr_27;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered5_wrport_we)
		storage_12[main_rtio_core_outputs_asyncfifobuffered5_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
	memadr_26 <= main_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_27 <= main_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r = storage_12[memadr_26];
assign main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r = storage_12[memadr_27];

reg [115:0] storage_13[0:127];
reg [6:0] memadr_28;
reg [6:0] memadr_29;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered6_wrport_we)
		storage_13[main_rtio_core_outputs_asyncfifobuffered6_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
	memadr_28 <= main_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_29 <= main_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r = storage_13[memadr_28];
assign main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r = storage_13[memadr_29];

reg [115:0] storage_14[0:127];
reg [6:0] memadr_30;
reg [6:0] memadr_31;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered7_wrport_we)
		storage_14[main_rtio_core_outputs_asyncfifobuffered7_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
	memadr_30 <= main_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_31 <= main_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r = storage_14[memadr_30];
assign main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r = storage_14[memadr_31];

reg [0:0] en_replaces_rom[0:36];
reg [5:0] memadr_32;
always @(posedge rio_clk) begin
	memadr_32 <= main_rtio_core_outputs_memory0_adr;
end

assign main_rtio_core_outputs_memory0_dat_r = en_replaces_rom[memadr_32];

initial begin
	$readmemh("en_replaces_rom.init", en_replaces_rom);
end

reg [0:0] en_replaces_rom_1[0:36];
reg [5:0] memadr_33;
always @(posedge rio_clk) begin
	memadr_33 <= main_rtio_core_outputs_memory1_adr;
end

assign main_rtio_core_outputs_memory1_dat_r = en_replaces_rom_1[memadr_33];

initial begin
	$readmemh("en_replaces_rom_1.init", en_replaces_rom_1);
end

reg [0:0] en_replaces_rom_2[0:36];
reg [5:0] memadr_34;
always @(posedge rio_clk) begin
	memadr_34 <= main_rtio_core_outputs_memory2_adr;
end

assign main_rtio_core_outputs_memory2_dat_r = en_replaces_rom_2[memadr_34];

initial begin
	$readmemh("en_replaces_rom_2.init", en_replaces_rom_2);
end

reg [0:0] en_replaces_rom_3[0:36];
reg [5:0] memadr_35;
always @(posedge rio_clk) begin
	memadr_35 <= main_rtio_core_outputs_memory3_adr;
end

assign main_rtio_core_outputs_memory3_dat_r = en_replaces_rom_3[memadr_35];

initial begin
	$readmemh("en_replaces_rom_3.init", en_replaces_rom_3);
end

reg [0:0] en_replaces_rom_4[0:36];
reg [5:0] memadr_36;
always @(posedge rio_clk) begin
	memadr_36 <= main_rtio_core_outputs_memory4_adr;
end

assign main_rtio_core_outputs_memory4_dat_r = en_replaces_rom_4[memadr_36];

initial begin
	$readmemh("en_replaces_rom_4.init", en_replaces_rom_4);
end

reg [0:0] en_replaces_rom_5[0:36];
reg [5:0] memadr_37;
always @(posedge rio_clk) begin
	memadr_37 <= main_rtio_core_outputs_memory5_adr;
end

assign main_rtio_core_outputs_memory5_dat_r = en_replaces_rom_5[memadr_37];

initial begin
	$readmemh("en_replaces_rom_5.init", en_replaces_rom_5);
end

reg [0:0] en_replaces_rom_6[0:36];
reg [5:0] memadr_38;
always @(posedge rio_clk) begin
	memadr_38 <= main_rtio_core_outputs_memory6_adr;
end

assign main_rtio_core_outputs_memory6_dat_r = en_replaces_rom_6[memadr_38];

initial begin
	$readmemh("en_replaces_rom_6.init", en_replaces_rom_6);
end

reg [0:0] en_replaces_rom_7[0:36];
reg [5:0] memadr_39;
always @(posedge rio_clk) begin
	memadr_39 <= main_rtio_core_outputs_memory7_adr;
end

assign main_rtio_core_outputs_memory7_dat_r = en_replaces_rom_7[memadr_39];

initial begin
	$readmemh("en_replaces_rom_7.init", en_replaces_rom_7);
end

reg [64:0] storage_15[0:63];
reg [5:0] memadr_40;
reg [5:0] memadr_41;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo0_wrport_we)
		storage_15[main_rtio_core_inputs_asyncfifo0_wrport_adr] <= main_rtio_core_inputs_asyncfifo0_wrport_dat_w;
	memadr_40 <= main_rtio_core_inputs_asyncfifo0_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_41 <= main_rtio_core_inputs_asyncfifo0_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo0_wrport_dat_r = storage_15[memadr_40];
assign main_rtio_core_inputs_asyncfifo0_rdport_dat_r = storage_15[memadr_41];

reg [64:0] storage_16[0:63];
reg [5:0] memadr_42;
reg [5:0] memadr_43;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo1_wrport_we)
		storage_16[main_rtio_core_inputs_asyncfifo1_wrport_adr] <= main_rtio_core_inputs_asyncfifo1_wrport_dat_w;
	memadr_42 <= main_rtio_core_inputs_asyncfifo1_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_43 <= main_rtio_core_inputs_asyncfifo1_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo1_wrport_dat_r = storage_16[memadr_42];
assign main_rtio_core_inputs_asyncfifo1_rdport_dat_r = storage_16[memadr_43];

reg [64:0] storage_17[0:63];
reg [5:0] memadr_44;
reg [5:0] memadr_45;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo2_wrport_we)
		storage_17[main_rtio_core_inputs_asyncfifo2_wrport_adr] <= main_rtio_core_inputs_asyncfifo2_wrport_dat_w;
	memadr_44 <= main_rtio_core_inputs_asyncfifo2_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_45 <= main_rtio_core_inputs_asyncfifo2_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo2_wrport_dat_r = storage_17[memadr_44];
assign main_rtio_core_inputs_asyncfifo2_rdport_dat_r = storage_17[memadr_45];

reg [64:0] storage_18[0:63];
reg [5:0] memadr_46;
reg [5:0] memadr_47;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo3_wrport_we)
		storage_18[main_rtio_core_inputs_asyncfifo3_wrport_adr] <= main_rtio_core_inputs_asyncfifo3_wrport_dat_w;
	memadr_46 <= main_rtio_core_inputs_asyncfifo3_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_47 <= main_rtio_core_inputs_asyncfifo3_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo3_wrport_dat_r = storage_18[memadr_46];
assign main_rtio_core_inputs_asyncfifo3_rdport_dat_r = storage_18[memadr_47];

reg [64:0] storage_19[0:63];
reg [5:0] memadr_48;
reg [5:0] memadr_49;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo4_wrport_we)
		storage_19[main_rtio_core_inputs_asyncfifo4_wrport_adr] <= main_rtio_core_inputs_asyncfifo4_wrport_dat_w;
	memadr_48 <= main_rtio_core_inputs_asyncfifo4_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_49 <= main_rtio_core_inputs_asyncfifo4_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo4_wrport_dat_r = storage_19[memadr_48];
assign main_rtio_core_inputs_asyncfifo4_rdport_dat_r = storage_19[memadr_49];

reg [64:0] storage_20[0:63];
reg [5:0] memadr_50;
reg [5:0] memadr_51;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo5_wrport_we)
		storage_20[main_rtio_core_inputs_asyncfifo5_wrport_adr] <= main_rtio_core_inputs_asyncfifo5_wrport_dat_w;
	memadr_50 <= main_rtio_core_inputs_asyncfifo5_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_51 <= main_rtio_core_inputs_asyncfifo5_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo5_wrport_dat_r = storage_20[memadr_50];
assign main_rtio_core_inputs_asyncfifo5_rdport_dat_r = storage_20[memadr_51];

reg [64:0] storage_21[0:63];
reg [5:0] memadr_52;
reg [5:0] memadr_53;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo6_wrport_we)
		storage_21[main_rtio_core_inputs_asyncfifo6_wrport_adr] <= main_rtio_core_inputs_asyncfifo6_wrport_dat_w;
	memadr_52 <= main_rtio_core_inputs_asyncfifo6_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_53 <= main_rtio_core_inputs_asyncfifo6_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo6_wrport_dat_r = storage_21[memadr_52];
assign main_rtio_core_inputs_asyncfifo6_rdport_dat_r = storage_21[memadr_53];

reg [64:0] storage_22[0:63];
reg [5:0] memadr_54;
reg [5:0] memadr_55;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo7_wrport_we)
		storage_22[main_rtio_core_inputs_asyncfifo7_wrport_adr] <= main_rtio_core_inputs_asyncfifo7_wrport_dat_w;
	memadr_54 <= main_rtio_core_inputs_asyncfifo7_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_55 <= main_rtio_core_inputs_asyncfifo7_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo7_wrport_dat_r = storage_22[memadr_54];
assign main_rtio_core_inputs_asyncfifo7_rdport_dat_r = storage_22[memadr_55];

reg [31:0] storage_23[0:3];
reg [1:0] memadr_56;
reg [1:0] memadr_57;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo8_wrport_we)
		storage_23[main_rtio_core_inputs_asyncfifo8_wrport_adr] <= main_rtio_core_inputs_asyncfifo8_wrport_dat_w;
	memadr_56 <= main_rtio_core_inputs_asyncfifo8_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_57 <= main_rtio_core_inputs_asyncfifo8_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo8_wrport_dat_r = storage_23[memadr_56];
assign main_rtio_core_inputs_asyncfifo8_rdport_dat_r = storage_23[memadr_57];

reg [31:0] storage_24[0:3];
reg [1:0] memadr_58;
reg [1:0] memadr_59;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo9_wrport_we)
		storage_24[main_rtio_core_inputs_asyncfifo9_wrport_adr] <= main_rtio_core_inputs_asyncfifo9_wrport_dat_w;
	memadr_58 <= main_rtio_core_inputs_asyncfifo9_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_59 <= main_rtio_core_inputs_asyncfifo9_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo9_wrport_dat_r = storage_24[memadr_58];
assign main_rtio_core_inputs_asyncfifo9_rdport_dat_r = storage_24[memadr_59];

reg [31:0] storage_25[0:3];
reg [1:0] memadr_60;
reg [1:0] memadr_61;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo10_wrport_we)
		storage_25[main_rtio_core_inputs_asyncfifo10_wrport_adr] <= main_rtio_core_inputs_asyncfifo10_wrport_dat_w;
	memadr_60 <= main_rtio_core_inputs_asyncfifo10_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_61 <= main_rtio_core_inputs_asyncfifo10_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo10_wrport_dat_r = storage_25[memadr_60];
assign main_rtio_core_inputs_asyncfifo10_rdport_dat_r = storage_25[memadr_61];

reg [256:0] storage_26[0:127];
reg [256:0] memdat_5;
reg [256:0] memdat_6;
always @(posedge sys_clk) begin
	if (main_rtio_analyzer_fifo_wrport_we)
		storage_26[main_rtio_analyzer_fifo_wrport_adr] <= main_rtio_analyzer_fifo_wrport_dat_w;
	memdat_5 <= storage_26[main_rtio_analyzer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (main_rtio_analyzer_fifo_rdport_re)
		memdat_6 <= storage_26[main_rtio_analyzer_fifo_rdport_adr];
end

assign main_rtio_analyzer_fifo_wrport_dat_r = memdat_5;
assign main_rtio_analyzer_fifo_rdport_dat_r = memdat_6;

reg [7:0] data_mem_grain0[0:8191];
reg [12:0] memadr_62;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[0])
		data_mem_grain0[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[7:0];
	memadr_62 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[7:0] = data_mem_grain0[memadr_62];

reg [7:0] data_mem_grain1[0:8191];
reg [12:0] memadr_63;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[1])
		data_mem_grain1[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[15:8];
	memadr_63 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[15:8] = data_mem_grain1[memadr_63];

reg [7:0] data_mem_grain2[0:8191];
reg [12:0] memadr_64;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[2])
		data_mem_grain2[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[23:16];
	memadr_64 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[23:16] = data_mem_grain2[memadr_64];

reg [7:0] data_mem_grain3[0:8191];
reg [12:0] memadr_65;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[3])
		data_mem_grain3[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[31:24];
	memadr_65 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[31:24] = data_mem_grain3[memadr_65];

reg [7:0] data_mem_grain4[0:8191];
reg [12:0] memadr_66;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[4])
		data_mem_grain4[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[39:32];
	memadr_66 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[39:32] = data_mem_grain4[memadr_66];

reg [7:0] data_mem_grain5[0:8191];
reg [12:0] memadr_67;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[5])
		data_mem_grain5[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[47:40];
	memadr_67 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[47:40] = data_mem_grain5[memadr_67];

reg [7:0] data_mem_grain6[0:8191];
reg [12:0] memadr_68;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[6])
		data_mem_grain6[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[55:48];
	memadr_68 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[55:48] = data_mem_grain6[memadr_68];

reg [7:0] data_mem_grain7[0:8191];
reg [12:0] memadr_69;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[7])
		data_mem_grain7[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[63:56];
	memadr_69 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[63:56] = data_mem_grain7[memadr_69];

reg [7:0] data_mem_grain8[0:8191];
reg [12:0] memadr_70;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[8])
		data_mem_grain8[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[71:64];
	memadr_70 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[71:64] = data_mem_grain8[memadr_70];

reg [7:0] data_mem_grain9[0:8191];
reg [12:0] memadr_71;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[9])
		data_mem_grain9[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[79:72];
	memadr_71 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[79:72] = data_mem_grain9[memadr_71];

reg [7:0] data_mem_grain10[0:8191];
reg [12:0] memadr_72;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[10])
		data_mem_grain10[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[87:80];
	memadr_72 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[87:80] = data_mem_grain10[memadr_72];

reg [7:0] data_mem_grain11[0:8191];
reg [12:0] memadr_73;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[11])
		data_mem_grain11[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[95:88];
	memadr_73 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[95:88] = data_mem_grain11[memadr_73];

reg [7:0] data_mem_grain12[0:8191];
reg [12:0] memadr_74;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[12])
		data_mem_grain12[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[103:96];
	memadr_74 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[103:96] = data_mem_grain12[memadr_74];

reg [7:0] data_mem_grain13[0:8191];
reg [12:0] memadr_75;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[13])
		data_mem_grain13[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[111:104];
	memadr_75 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[111:104] = data_mem_grain13[memadr_75];

reg [7:0] data_mem_grain14[0:8191];
reg [12:0] memadr_76;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[14])
		data_mem_grain14[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[119:112];
	memadr_76 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[119:112] = data_mem_grain14[memadr_76];

reg [7:0] data_mem_grain15[0:8191];
reg [12:0] memadr_77;
always @(posedge sys_clk) begin
	if (main_genericstandalone_genericstandalone_genericstandalone_data_port_we[15])
		data_mem_grain15[main_genericstandalone_genericstandalone_genericstandalone_data_port_adr] <= main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_w[127:120];
	memadr_77 <= main_genericstandalone_genericstandalone_genericstandalone_data_port_adr;
end

assign main_genericstandalone_genericstandalone_genericstandalone_data_port_dat_r[127:120] = data_mem_grain15[memadr_77];

reg [7:0] mem_grain0[0:381];
reg [8:0] memadr_78;
reg [8:0] memadr_79;
always @(posedge sys_clk) begin
	memadr_78 <= main_genericstandalone_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram0_we[0])
		mem_grain0[main_genericstandalone_sram0_adr1] <= main_genericstandalone_sram0_dat_w[7:0];
	memadr_79 <= main_genericstandalone_sram0_adr1;
end

assign main_genericstandalone_reader_memory0_dat_r[7:0] = mem_grain0[memadr_78];
assign main_genericstandalone_sram0_dat_r1[7:0] = mem_grain0[memadr_79];

reg [7:0] mem_grain1[0:381];
reg [8:0] memadr_80;
reg [8:0] memadr_81;
always @(posedge sys_clk) begin
	memadr_80 <= main_genericstandalone_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram0_we[1])
		mem_grain1[main_genericstandalone_sram0_adr1] <= main_genericstandalone_sram0_dat_w[15:8];
	memadr_81 <= main_genericstandalone_sram0_adr1;
end

assign main_genericstandalone_reader_memory0_dat_r[15:8] = mem_grain1[memadr_80];
assign main_genericstandalone_sram0_dat_r1[15:8] = mem_grain1[memadr_81];

reg [7:0] mem_grain2[0:381];
reg [8:0] memadr_82;
reg [8:0] memadr_83;
always @(posedge sys_clk) begin
	memadr_82 <= main_genericstandalone_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram0_we[2])
		mem_grain2[main_genericstandalone_sram0_adr1] <= main_genericstandalone_sram0_dat_w[23:16];
	memadr_83 <= main_genericstandalone_sram0_adr1;
end

assign main_genericstandalone_reader_memory0_dat_r[23:16] = mem_grain2[memadr_82];
assign main_genericstandalone_sram0_dat_r1[23:16] = mem_grain2[memadr_83];

reg [7:0] mem_grain3[0:381];
reg [8:0] memadr_84;
reg [8:0] memadr_85;
always @(posedge sys_clk) begin
	memadr_84 <= main_genericstandalone_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram0_we[3])
		mem_grain3[main_genericstandalone_sram0_adr1] <= main_genericstandalone_sram0_dat_w[31:24];
	memadr_85 <= main_genericstandalone_sram0_adr1;
end

assign main_genericstandalone_reader_memory0_dat_r[31:24] = mem_grain3[memadr_84];
assign main_genericstandalone_sram0_dat_r1[31:24] = mem_grain3[memadr_85];

reg [7:0] mem_grain0_1[0:381];
reg [8:0] memadr_86;
reg [8:0] memadr_87;
always @(posedge sys_clk) begin
	memadr_86 <= main_genericstandalone_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram1_we[0])
		mem_grain0_1[main_genericstandalone_sram1_adr1] <= main_genericstandalone_sram1_dat_w[7:0];
	memadr_87 <= main_genericstandalone_sram1_adr1;
end

assign main_genericstandalone_reader_memory1_dat_r[7:0] = mem_grain0_1[memadr_86];
assign main_genericstandalone_sram1_dat_r1[7:0] = mem_grain0_1[memadr_87];

reg [7:0] mem_grain1_1[0:381];
reg [8:0] memadr_88;
reg [8:0] memadr_89;
always @(posedge sys_clk) begin
	memadr_88 <= main_genericstandalone_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram1_we[1])
		mem_grain1_1[main_genericstandalone_sram1_adr1] <= main_genericstandalone_sram1_dat_w[15:8];
	memadr_89 <= main_genericstandalone_sram1_adr1;
end

assign main_genericstandalone_reader_memory1_dat_r[15:8] = mem_grain1_1[memadr_88];
assign main_genericstandalone_sram1_dat_r1[15:8] = mem_grain1_1[memadr_89];

reg [7:0] mem_grain2_1[0:381];
reg [8:0] memadr_90;
reg [8:0] memadr_91;
always @(posedge sys_clk) begin
	memadr_90 <= main_genericstandalone_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram1_we[2])
		mem_grain2_1[main_genericstandalone_sram1_adr1] <= main_genericstandalone_sram1_dat_w[23:16];
	memadr_91 <= main_genericstandalone_sram1_adr1;
end

assign main_genericstandalone_reader_memory1_dat_r[23:16] = mem_grain2_1[memadr_90];
assign main_genericstandalone_sram1_dat_r1[23:16] = mem_grain2_1[memadr_91];

reg [7:0] mem_grain3_1[0:381];
reg [8:0] memadr_92;
reg [8:0] memadr_93;
always @(posedge sys_clk) begin
	memadr_92 <= main_genericstandalone_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram1_we[3])
		mem_grain3_1[main_genericstandalone_sram1_adr1] <= main_genericstandalone_sram1_dat_w[31:24];
	memadr_93 <= main_genericstandalone_sram1_adr1;
end

assign main_genericstandalone_reader_memory1_dat_r[31:24] = mem_grain3_1[memadr_92];
assign main_genericstandalone_sram1_dat_r1[31:24] = mem_grain3_1[memadr_93];

reg [7:0] mem_grain0_2[0:381];
reg [8:0] memadr_94;
reg [8:0] memadr_95;
always @(posedge sys_clk) begin
	memadr_94 <= main_genericstandalone_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram2_we[0])
		mem_grain0_2[main_genericstandalone_sram2_adr1] <= main_genericstandalone_sram2_dat_w[7:0];
	memadr_95 <= main_genericstandalone_sram2_adr1;
end

assign main_genericstandalone_reader_memory2_dat_r[7:0] = mem_grain0_2[memadr_94];
assign main_genericstandalone_sram2_dat_r1[7:0] = mem_grain0_2[memadr_95];

reg [7:0] mem_grain1_2[0:381];
reg [8:0] memadr_96;
reg [8:0] memadr_97;
always @(posedge sys_clk) begin
	memadr_96 <= main_genericstandalone_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram2_we[1])
		mem_grain1_2[main_genericstandalone_sram2_adr1] <= main_genericstandalone_sram2_dat_w[15:8];
	memadr_97 <= main_genericstandalone_sram2_adr1;
end

assign main_genericstandalone_reader_memory2_dat_r[15:8] = mem_grain1_2[memadr_96];
assign main_genericstandalone_sram2_dat_r1[15:8] = mem_grain1_2[memadr_97];

reg [7:0] mem_grain2_2[0:381];
reg [8:0] memadr_98;
reg [8:0] memadr_99;
always @(posedge sys_clk) begin
	memadr_98 <= main_genericstandalone_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram2_we[2])
		mem_grain2_2[main_genericstandalone_sram2_adr1] <= main_genericstandalone_sram2_dat_w[23:16];
	memadr_99 <= main_genericstandalone_sram2_adr1;
end

assign main_genericstandalone_reader_memory2_dat_r[23:16] = mem_grain2_2[memadr_98];
assign main_genericstandalone_sram2_dat_r1[23:16] = mem_grain2_2[memadr_99];

reg [7:0] mem_grain3_2[0:381];
reg [8:0] memadr_100;
reg [8:0] memadr_101;
always @(posedge sys_clk) begin
	memadr_100 <= main_genericstandalone_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram2_we[3])
		mem_grain3_2[main_genericstandalone_sram2_adr1] <= main_genericstandalone_sram2_dat_w[31:24];
	memadr_101 <= main_genericstandalone_sram2_adr1;
end

assign main_genericstandalone_reader_memory2_dat_r[31:24] = mem_grain3_2[memadr_100];
assign main_genericstandalone_sram2_dat_r1[31:24] = mem_grain3_2[memadr_101];

reg [7:0] mem_grain0_3[0:381];
reg [8:0] memadr_102;
reg [8:0] memadr_103;
always @(posedge sys_clk) begin
	memadr_102 <= main_genericstandalone_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram3_we[0])
		mem_grain0_3[main_genericstandalone_sram3_adr1] <= main_genericstandalone_sram3_dat_w[7:0];
	memadr_103 <= main_genericstandalone_sram3_adr1;
end

assign main_genericstandalone_reader_memory3_dat_r[7:0] = mem_grain0_3[memadr_102];
assign main_genericstandalone_sram3_dat_r1[7:0] = mem_grain0_3[memadr_103];

reg [7:0] mem_grain1_3[0:381];
reg [8:0] memadr_104;
reg [8:0] memadr_105;
always @(posedge sys_clk) begin
	memadr_104 <= main_genericstandalone_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram3_we[1])
		mem_grain1_3[main_genericstandalone_sram3_adr1] <= main_genericstandalone_sram3_dat_w[15:8];
	memadr_105 <= main_genericstandalone_sram3_adr1;
end

assign main_genericstandalone_reader_memory3_dat_r[15:8] = mem_grain1_3[memadr_104];
assign main_genericstandalone_sram3_dat_r1[15:8] = mem_grain1_3[memadr_105];

reg [7:0] mem_grain2_3[0:381];
reg [8:0] memadr_106;
reg [8:0] memadr_107;
always @(posedge sys_clk) begin
	memadr_106 <= main_genericstandalone_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram3_we[2])
		mem_grain2_3[main_genericstandalone_sram3_adr1] <= main_genericstandalone_sram3_dat_w[23:16];
	memadr_107 <= main_genericstandalone_sram3_adr1;
end

assign main_genericstandalone_reader_memory3_dat_r[23:16] = mem_grain2_3[memadr_106];
assign main_genericstandalone_sram3_dat_r1[23:16] = mem_grain2_3[memadr_107];

reg [7:0] mem_grain3_3[0:381];
reg [8:0] memadr_108;
reg [8:0] memadr_109;
always @(posedge sys_clk) begin
	memadr_108 <= main_genericstandalone_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_genericstandalone_sram3_we[3])
		mem_grain3_3[main_genericstandalone_sram3_adr1] <= main_genericstandalone_sram3_dat_w[31:24];
	memadr_109 <= main_genericstandalone_sram3_adr1;
end

assign main_genericstandalone_reader_memory3_dat_r[31:24] = mem_grain3_3[memadr_108];
assign main_genericstandalone_sram3_dat_r1[31:24] = mem_grain3_3[memadr_109];

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(builder_xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(clk200_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(builder_xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(eth_tx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2),
	.Q(builder_xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2),
	.Q(eth_rx_rst)
);

OBUFDS OBUFDS_1(
	.I(main_pad0),
	.O(urukul2_dds_reset_sync_in_p),
	.OB(urukul2_dds_reset_sync_in_n)
);

OBUFDS OBUFDS_2(
	.I(main_pad1),
	.O(urukul4_dds_reset_sync_in_p),
	.OB(urukul4_dds_reset_sync_in_n)
);

OBUFDS OBUFDS_3(
	.I(main_pad2),
	.O(urukul6_dds_reset_sync_in_p),
	.OB(urukul6_dds_reset_sync_in_n)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl3),
	.Q(builder_xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl3),
	.Q(rtio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(rio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_rtio_core_cmd_reset),
	.Q(builder_xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(rio_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(main_rtio_core_cmd_reset),
	.Q(rio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_rtio_core_cmd_reset_phy),
	.Q(builder_xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(main_rtio_core_cmd_reset_phy),
	.Q(rio_phy_rst)
);

endmodule
