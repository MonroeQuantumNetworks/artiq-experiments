/* Machine-generated using Migen */
module top(
	input serial_rx,
	output reg serial_tx,
	input clk125_gtp_p,
	input clk125_gtp_n,
	output [14:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash2x_cs_n,
	inout [1:0] spiflash2x_dq,
	input spiflash2x_wp,
	input spiflash2x_hold,
	output sfp_txp,
	output sfp_txn,
	input sfp_rxp,
	input sfp_rxn,
	input sfp_ctl_mod_def1,
	input sfp_ctl_mod_def2,
	input sfp_ctl_los,
	input sfp_ctl_mod_present,
	output sfp_ctl_rate_select,
	output sfp_ctl_tx_disable,
	input sfp_ctl_tx_fault,
	output sfp_ctl_led,
	output user_led,
	inout i2c_scl,
	inout i2c_sda,
	output clk_sel,
	inout dio0_p,
	inout dio0_n,
	inout dio0_p_1,
	inout dio0_n_1,
	inout dio0_p_2,
	inout dio0_n_2,
	inout dio0_p_3,
	inout dio0_n_3,
	inout dio0_p_4,
	inout dio0_n_4,
	inout dio0_p_5,
	inout dio0_n_5,
	inout dio0_p_6,
	inout dio0_n_6,
	inout dio0_p_7,
	inout dio0_n_7,
	inout dio1_p,
	inout dio1_n,
	inout dio1_p_1,
	inout dio1_n_1,
	inout dio1_p_2,
	inout dio1_n_2,
	inout dio1_p_3,
	inout dio1_n_3,
	inout dio1_p_4,
	inout dio1_n_4,
	inout dio1_p_5,
	inout dio1_n_5,
	inout dio1_p_6,
	inout dio1_n_6,
	inout dio1_p_7,
	inout dio1_n_7,
	output urukul2_spi_p_clk,
	inout urukul2_spi_p_mosi,
	inout urukul2_spi_p_miso,
	output [2:0] urukul2_spi_p_cs_n,
	output urukul2_spi_n_clk,
	inout urukul2_spi_n_mosi,
	inout urukul2_spi_n_miso,
	output [2:0] urukul2_spi_n_cs_n,
	output urukul2_dds_reset_sync_in_p,
	output urukul2_dds_reset_sync_in_n,
	inout urukul2_io_update_p,
	inout urukul2_io_update_n,
	inout urukul2_sw0_p,
	inout urukul2_sw0_n,
	inout urukul2_sw1_p,
	inout urukul2_sw1_n,
	inout urukul2_sw2_p,
	inout urukul2_sw2_n,
	inout urukul2_sw3_p,
	inout urukul2_sw3_n,
	output urukul4_spi_p_clk,
	inout urukul4_spi_p_mosi,
	inout urukul4_spi_p_miso,
	output [2:0] urukul4_spi_p_cs_n,
	output urukul4_spi_n_clk,
	inout urukul4_spi_n_mosi,
	inout urukul4_spi_n_miso,
	output [2:0] urukul4_spi_n_cs_n,
	output urukul4_dds_reset_sync_in_p,
	output urukul4_dds_reset_sync_in_n,
	inout urukul4_io_update_p,
	inout urukul4_io_update_n,
	inout urukul4_sw0_p,
	inout urukul4_sw0_n,
	inout urukul4_sw1_p,
	inout urukul4_sw1_n,
	inout urukul4_sw2_p,
	inout urukul4_sw2_n,
	inout urukul4_sw3_p,
	inout urukul4_sw3_n,
	output urukul6_spi_p_clk,
	inout urukul6_spi_p_mosi,
	inout urukul6_spi_p_miso,
	output [2:0] urukul6_spi_p_cs_n,
	output urukul6_spi_n_clk,
	inout urukul6_spi_n_mosi,
	inout urukul6_spi_n_miso,
	output [2:0] urukul6_spi_n_cs_n,
	output urukul6_dds_reset_sync_in_p,
	output urukul6_dds_reset_sync_in_n,
	inout urukul6_io_update_p,
	inout urukul6_io_update_n,
	inout urukul6_sw0_p,
	inout urukul6_sw0_n,
	inout urukul6_sw1_p,
	inout urukul6_sw1_n,
	inout urukul6_sw2_p,
	inout urukul6_sw2_n,
	inout urukul6_sw3_p,
	inout urukul6_sw3_n,
	input sfp_ctl_mod_def1_1,
	input sfp_ctl_mod_def2_1,
	input sfp_ctl_los_1,
	input sfp_ctl_mod_present_1,
	input sfp_ctl_rate_select_1,
	input sfp_ctl_tx_disable_1,
	input sfp_ctl_tx_fault_1,
	output sfp_ctl_led_1,
	input sfp_ctl_mod_def1_2,
	input sfp_ctl_mod_def2_2,
	input sfp_ctl_los_2,
	input sfp_ctl_mod_present_2,
	input sfp_ctl_rate_select_2,
	input sfp_ctl_tx_disable_2,
	input sfp_ctl_tx_fault_2,
	output sfp_ctl_led_2,
	input si5324_clkout_fabric_p,
	input si5324_clkout_fabric_n
);

wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_bte;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_err;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_err;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_i_adr_o;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_d_adr_o;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_bte;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_err;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_re = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_re = 1'd0;
reg [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full = 30'd0;
wire [17:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_re = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error = 1'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_err = 1'd0;
wire [9:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_r;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w;
reg [13:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr = 14'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we = 1'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w = 8'd0;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_r;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_err = 1'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter = 2'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full = 32'd4367715;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_payload_data;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg = 8'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount = 4'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_stb = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_ack;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_eop = 1'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_payload_data = 8'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_rx = 32'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_r = 1'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_reg = 8'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount = 4'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_re;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_r;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_w;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_txfull_status;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxempty_status;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_irq;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_status;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_pending = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_trigger;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_clear;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_old_trigger = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_status;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_pending = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_trigger;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_clear;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_old_trigger = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_re;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_r;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_w;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_re;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_r;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_ack;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_eop = 1'd0;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_readable;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_din;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_dout;
reg [4:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level = 5'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_replace = 1'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce = 4'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_consume = 4'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_we;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_dat_w;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_do_read;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_adr;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_dat_r;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_eop;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_readable;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_din;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_dout;
reg [4:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level = 5'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_replace = 1'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce = 4'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_consume = 4'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_we;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_dat_w;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_do_read;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_adr;
wire [8:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_dat_r;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_payload_data;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_eop;
reg [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full = 64'd0;
wire [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_re = 1'd0;
reg [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full = 64'd0;
wire [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_re = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_w = 1'd0;
reg [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status = 64'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_irq;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_status;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_pending = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_trigger;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_clear;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_old_trigger = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_r;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_w;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_r;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_w;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_re = 1'd0;
reg [63:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value = 64'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_buf;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_div2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_locked;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_fb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x_dqs;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_locked;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_fb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_clk200;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_meta;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_unbuf;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_reset_counter = 4'd15;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ic_reset = 1'd1;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_w = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_w = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_sd_clk_se;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dqs = 1'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern = 8'd85;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t1;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o8;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay8;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed8;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t8;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o9;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay9;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed9;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t9;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o10;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay10;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed10;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t10;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o11;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay11;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed11;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t11;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o12;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay12;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed12;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t12;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o13;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay13;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed13;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t13;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o14;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay14;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed14;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t14;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o15;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay15;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed15;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t15;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en0 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en1 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en2 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en3 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en = 4'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_bte;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_err;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_valid;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_bank;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cs_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_ras_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_mask;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_en;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_address;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_we_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cke;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_odt;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_reset_n;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_en;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_address;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_we_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cke;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_odt;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_reset_n;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_en;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_address;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_we_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cke;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_odt;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_reset_n;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_en;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_address;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cas_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_we_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cke;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_odt;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_reset_n;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_en;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_valid;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage_full = 4'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_re = 1'd0;
reg [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_w = 1'd0;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full = 15'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_re = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status = 32'd0;
reg [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_w = 1'd0;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full = 15'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_re = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status = 32'd0;
reg [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_w = 1'd0;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full = 15'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_re = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full = 32'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status = 32'd0;
reg [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_re;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_w = 1'd0;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full = 15'd0;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_re = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full = 32'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status = 32'd0;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata_en = 1'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata_en = 1'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata_en = 1'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_en;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cas_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_ras_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_we_n;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_en;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata_en = 1'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata_valid;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_bank;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cas_n = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cs_n;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_ras_n = 1'd1;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_we_n = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cke;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_odt;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_reset_n;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata_en = 1'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata_mask;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata_en = 1'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata_valid;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr;
wire [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_w;
wire [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_r;
wire [15:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_err = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_idle;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_hit;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset2;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset3;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset5;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset6;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_open;
wire [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_hit;
reg [14:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row1 = 15'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset7;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_wait;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_done;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count = 3'd4;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_wait;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_done;
reg [9:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count = 10'd886;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_adr;
wire [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_w;
wire [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_r;
wire [15:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_sel;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_stb;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_ack;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_we;
reg [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cti = 3'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_bte = 2'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_err;
wire [12:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
wire [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r;
reg [15:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we;
reg [127:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_write_from_slave;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_adr_offset_r = 2'd0;
wire [12:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_adr;
wire [19:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_r;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_we;
wire [19:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_w;
wire [18:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_tag;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_dirty;
wire [18:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_tag;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_dirty;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_clr;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_inc;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk;
wire [29:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_err = 1'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage_full = 4'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_re = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_status;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_re = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_cs_n = 1'd1;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_clk = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dq_oe = 1'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_o;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe;
wire [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr = 32'd0;
reg monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 = 1'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dqi = 2'd0;
reg [6:0] monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter = 7'd0;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_reset;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_lock;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_clk;
wire monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_refclk;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb;
wire [15:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg;
wire monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_stb;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_ack;
wire [7:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_data;
reg [7:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0;
reg [9:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output0 = 10'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disparity = 1'd0;
wire [7:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1;
wire monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k1;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_in = 1'd0;
reg [9:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out;
reg [5:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b = 6'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_unbalanced = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_flip = 1'd0;
reg [3:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b = 4'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_unbalanced = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_flip = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1 = 1'd0;
reg [5:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_6b;
wire monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter;
reg [3:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b;
wire [9:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_parity = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type = 1'd0;
reg [15:0] monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg_buffer = 16'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_load_config_reg_buffer;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en;
wire [7:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_data;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_valid_ci;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg = 1'd0;
reg [15:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg = 16'd0;
wire [9:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input;
wire [7:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k = 1'd0;
reg [9:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first;
reg [4:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code5b = 5'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b = 3'd0;
reg [7:0] monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg_lsb = 8'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_lsb;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_msb;
reg monroe_ionphoton_monroe_ionphoton_pcs_receivepath_first_preamble_byte;
wire monroe_ionphoton_monroe_ionphoton_pcs_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_pcs_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_pcs_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_pcs_source_stb = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_source_ack;
wire monroe_ionphoton_monroe_ionphoton_pcs_source_eop;
reg [7:0] monroe_ionphoton_monroe_ionphoton_pcs_source_payload_data = 8'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_source_payload_last_be = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_source_payload_error = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_link_up;
reg monroe_ionphoton_monroe_ionphoton_pcs_restart;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_en_d = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_i;
wire monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o_r = 1'd0;
reg [19:0] monroe_ionphoton_monroe_ionphoton_pcs_checker_counter = 20'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_checker_tick = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_checker_ok = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_autoneg_ack;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o_r = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_pcs_wait;
wire monroe_ionphoton_monroe_ionphoton_pcs_done;
reg [20:0] monroe_ionphoton_monroe_ionphoton_pcs_count = 21'd1250000;
reg [2:0] monroe_ionphoton_monroe_ionphoton_pcs_c_counter = 3'd0;
reg [15:0] monroe_ionphoton_monroe_ionphoton_pcs_previous_config_reg = 16'd0;
wire eth_tx_clk;
wire eth_tx_rst;
wire eth_rx_clk;
wire eth_rx_rst;
wire eth_tx_half_clk;
wire eth_rx_half_clk;
wire monroe_ionphoton_monroe_ionphoton_txoutclk;
wire monroe_ionphoton_monroe_ionphoton_rxoutclk;
wire monroe_ionphoton_monroe_ionphoton_tx_reset;
wire monroe_ionphoton_monroe_ionphoton_tx_mmcm_locked;
wire [19:0] monroe_ionphoton_monroe_ionphoton_tx_data0;
wire monroe_ionphoton_monroe_ionphoton_tx_reset_done;
wire monroe_ionphoton_monroe_ionphoton_rx_reset;
wire monroe_ionphoton_monroe_ionphoton_rx_mmcm_locked;
wire [19:0] monroe_ionphoton_monroe_ionphoton_rx_data0;
wire monroe_ionphoton_monroe_ionphoton_rx_reset_done;
wire monroe_ionphoton_monroe_ionphoton_rx_pma_reset_done;
wire [8:0] monroe_ionphoton_monroe_ionphoton_drpaddr;
wire monroe_ionphoton_monroe_ionphoton_drpen;
wire [15:0] monroe_ionphoton_monroe_ionphoton_drpdi;
wire monroe_ionphoton_monroe_ionphoton_drprdy;
wire [15:0] monroe_ionphoton_monroe_ionphoton_drpdo;
wire monroe_ionphoton_monroe_ionphoton_drpwe;
wire monroe_ionphoton_monroe_ionphoton_txoutclk_rebuffer;
wire monroe_ionphoton_monroe_ionphoton_rxoutclk_rebuffer;
wire monroe_ionphoton_monroe_ionphoton_tx_mmcm_fb;
(* dont_touch = "true" *) reg monroe_ionphoton_monroe_ionphoton_tx_mmcm_reset = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_clk_tx_unbuf;
wire monroe_ionphoton_monroe_ionphoton_clk_tx_half_unbuf;
wire monroe_ionphoton_monroe_ionphoton_rx_mmcm_fb;
(* dont_touch = "true" *) reg monroe_ionphoton_monroe_ionphoton_rx_mmcm_reset = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_clk_rx_unbuf;
wire monroe_ionphoton_monroe_ionphoton_clk_rx_half_unbuf;
(* dont_touch = "true" *) reg monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock0;
(* dont_touch = "true" *) reg monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset0 = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_tx_init_done;
reg monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset1;
reg monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset1;
wire monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock1;
reg [5:0] monroe_ionphoton_monroe_ionphoton_tx_init_timer = 6'd0;
reg monroe_ionphoton_monroe_ionphoton_tx_init_tick = 1'd0;
(* dont_touch = "true" *) reg monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_rx_init_drpaddr;
reg monroe_ionphoton_monroe_ionphoton_rx_init_drpen;
reg [15:0] monroe_ionphoton_monroe_ionphoton_rx_init_drpdi;
wire monroe_ionphoton_monroe_ionphoton_rx_init_drprdy;
wire [15:0] monroe_ionphoton_monroe_ionphoton_rx_init_drpdo;
reg monroe_ionphoton_monroe_ionphoton_rx_init_drpwe;
wire monroe_ionphoton_monroe_ionphoton_rx_init_enable;
wire monroe_ionphoton_monroe_ionphoton_rx_init_restart;
reg monroe_ionphoton_monroe_ionphoton_rx_init_done;
reg monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1;
wire monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done1;
reg [15:0] monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue = 16'd0;
reg monroe_ionphoton_monroe_ionphoton_rx_init_drpmask;
reg monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done_r = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_i;
wire monroe_ionphoton_monroe_ionphoton_o;
reg monroe_ionphoton_monroe_ionphoton_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_toggle_o_r = 1'd0;
reg [12:0] monroe_ionphoton_monroe_ionphoton_cdr_lock_counter = 13'd0;
reg monroe_ionphoton_monroe_ionphoton_cdr_locked = 1'd0;
wire [9:0] monroe_ionphoton_monroe_ionphoton_tx_data1;
reg [19:0] monroe_ionphoton_monroe_ionphoton_tx_data_half = 20'd0;
wire [19:0] monroe_ionphoton_monroe_ionphoton_rx_data_half;
reg [9:0] monroe_ionphoton_monroe_ionphoton_rx_data1 = 10'd0;
reg [19:0] monroe_ionphoton_monroe_ionphoton_buf = 20'd0;
reg monroe_ionphoton_monroe_ionphoton_phase_half = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_phase_half_rereg = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_ack;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_eop;
reg [7:0] monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_data;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_error;
reg [3:0] monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter = 4'd0;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_reset;
reg monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_ce;
reg [31:0] monroe_ionphoton_monroe_ionphoton_preamble_errors_status = 32'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_crc_errors_status = 32'd0;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_eop;
reg [7:0] monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_error;
reg [63:0] monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt = 3'd0;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_clr_cnt;
reg monroe_ionphoton_monroe_ionphoton_preamble_inserter_inc_cnt;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_preamble_checker_source_stb;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_source_ack;
reg monroe_ionphoton_monroe_ionphoton_preamble_checker_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_error;
reg monroe_ionphoton_monroe_ionphoton_preamble_checker_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop;
reg [7:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_error;
reg [7:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_data0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_value;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_error;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_last;
reg [31:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_next;
reg [31:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg = 32'd4294967295;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_ce;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_reset;
reg [1:0] monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt = 2'd3;
wire monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt_done;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing0;
reg monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing1;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_stb;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_ack;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_error;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_value;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_error;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last;
reg [31:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next;
reg [31:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg = 32'd4294967295;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_ce;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reset;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_stb;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_ack;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_readable;
wire [10:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_din;
wire [10:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level = 3'd0;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr;
wire [10:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_we;
wire [10:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_dat_w;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_do_read;
wire [2:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_adr;
wire [10:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_data;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_error;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_eop;
reg monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_reset;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_in;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_out;
wire monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_full;
wire monroe_ionphoton_monroe_ionphoton_ps_preamble_error_i;
wire monroe_ionphoton_monroe_ionphoton_ps_preamble_error_o;
reg monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o_r = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_ps_crc_error_i;
wire monroe_ionphoton_monroe_ionphoton_ps_crc_error_o;
reg monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_i = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o;
reg monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o_r = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_error;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_source_ack;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop;
reg [7:0] monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_data;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_last_be;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_error;
reg [15:0] monroe_ionphoton_monroe_ionphoton_padding_inserter_counter = 16'd1;
wire monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_done;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_reset;
reg monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_ce;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_source_stb;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_source_ack;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_source_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_source_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_last_be_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_data;
reg monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_last_be = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_error = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_tx_last_be_ongoing = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_source_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_source_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_data;
reg monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_data;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_eop;
reg [39:0] monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_eop;
reg [9:0] monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data;
reg [1:0] monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux = 2'd0;
wire monroe_ionphoton_monroe_ionphoton_tx_converter_converter_last;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_eop;
wire [7:0] monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_last_be;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_eop;
reg [31:0] monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data;
reg [3:0] monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be;
reg [3:0] monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_eop;
wire [9:0] monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_ack;
reg monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop = 1'd0;
reg [39:0] monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data = 40'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux = 2'd0;
wire monroe_ionphoton_monroe_ionphoton_rx_converter_converter_load_part;
reg monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_source_stb;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_source_ack;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_source_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_readable;
wire [40:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_din;
wire [40:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_dout;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next;
reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next;
reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary;
wire [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_produce_rdomain;
wire [6:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_consume_wdomain;
wire [5:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_adr;
wire [40:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_we;
wire [40:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_dat_w;
wire [5:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_adr;
wire [40:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_dat_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_error;
wire monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_eop;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_source_stb;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_source_ack;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_source_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_readable;
wire [40:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_din;
wire [40:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_dout;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next;
reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next;
reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary;
wire [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_produce_rdomain;
wire [6:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_consume_wdomain;
wire [5:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_adr;
wire [40:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_we;
wire [40:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_dat_w;
wire [5:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_adr;
wire [40:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_dat_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_error;
wire monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_eop;
wire monroe_ionphoton_monroe_ionphoton_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_sink_ack;
wire monroe_ionphoton_monroe_ionphoton_sink_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sink_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sink_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sink_payload_error;
wire monroe_ionphoton_monroe_ionphoton_source_stb;
wire monroe_ionphoton_monroe_ionphoton_source_ack;
wire monroe_ionphoton_monroe_ionphoton_source_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_source_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_source_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_source_payload_error;
wire [29:0] monroe_ionphoton_monroe_ionphoton_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_bus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_bus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_bus_stb;
wire monroe_ionphoton_monroe_ionphoton_bus_ack;
wire monroe_ionphoton_monroe_ionphoton_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_bus_bte;
wire monroe_ionphoton_monroe_ionphoton_bus_err;
wire monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb;
reg monroe_ionphoton_monroe_ionphoton_writer_sink_sink_ack = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_writer_sink_sink_eop;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data;
wire [3:0] monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be;
wire [3:0] monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_error;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_slot_status;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_length_status;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_errors_status = 32'd0;
wire monroe_ionphoton_monroe_ionphoton_writer_irq;
wire monroe_ionphoton_monroe_ionphoton_writer_available_status;
wire monroe_ionphoton_monroe_ionphoton_writer_available_pending;
wire monroe_ionphoton_monroe_ionphoton_writer_available_trigger;
reg monroe_ionphoton_monroe_ionphoton_writer_available_clear;
wire monroe_ionphoton_monroe_ionphoton_writer_status_re;
wire monroe_ionphoton_monroe_ionphoton_writer_status_r;
wire monroe_ionphoton_monroe_ionphoton_writer_status_w;
wire monroe_ionphoton_monroe_ionphoton_writer_pending_re;
wire monroe_ionphoton_monroe_ionphoton_writer_pending_r;
wire monroe_ionphoton_monroe_ionphoton_writer_pending_w;
reg monroe_ionphoton_monroe_ionphoton_writer_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_writer_storage;
reg monroe_ionphoton_monroe_ionphoton_writer_re = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_writer_increment;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_counter = 32'd0;
reg monroe_ionphoton_monroe_ionphoton_writer_counter_reset;
reg monroe_ionphoton_monroe_ionphoton_writer_counter_ce;
reg [1:0] monroe_ionphoton_monroe_ionphoton_writer_slot = 2'd0;
reg monroe_ionphoton_monroe_ionphoton_writer_slot_ce;
reg monroe_ionphoton_monroe_ionphoton_writer_ongoing;
reg monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_ack;
reg monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_eop = 1'd0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_slot;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_length;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_source_stb;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_source_ack;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_source_eop;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_slot;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_length;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_readable;
wire [34:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_din;
wire [34:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_dout;
reg [2:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_level = 3'd0;
reg monroe_ionphoton_monroe_ionphoton_writer_fifo_replace = 1'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_produce = 2'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_consume = 2'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr;
wire [34:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_we;
wire [34:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_dat_w;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_do_read;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_adr;
wire [34:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_dat_r;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_slot;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_length;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_eop;
wire [1:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_slot;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_length;
wire monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_eop;
reg [8:0] monroe_ionphoton_monroe_ionphoton_writer_memory0_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_r;
reg monroe_ionphoton_monroe_ionphoton_writer_memory0_we;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_w;
reg [8:0] monroe_ionphoton_monroe_ionphoton_writer_memory1_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_r;
reg monroe_ionphoton_monroe_ionphoton_writer_memory1_we;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_w;
reg [8:0] monroe_ionphoton_monroe_ionphoton_writer_memory2_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_r;
reg monroe_ionphoton_monroe_ionphoton_writer_memory2_we;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_w;
reg [8:0] monroe_ionphoton_monroe_ionphoton_writer_memory3_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_r;
reg monroe_ionphoton_monroe_ionphoton_writer_memory3_we;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_w;
reg monroe_ionphoton_monroe_ionphoton_reader_source_source_stb;
wire monroe_ionphoton_monroe_ionphoton_reader_source_source_ack;
reg monroe_ionphoton_monroe_ionphoton_reader_source_source_eop;
reg [31:0] monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data;
reg [3:0] monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be;
reg [3:0] monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_error = 4'd0;
wire monroe_ionphoton_monroe_ionphoton_reader_start_re;
wire monroe_ionphoton_monroe_ionphoton_reader_start_r;
reg monroe_ionphoton_monroe_ionphoton_reader_start_w = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_reader_ready_status;
reg [1:0] monroe_ionphoton_monroe_ionphoton_reader_slot_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_slot_storage;
reg monroe_ionphoton_monroe_ionphoton_reader_slot_re = 1'd0;
reg [10:0] monroe_ionphoton_monroe_ionphoton_reader_length_storage_full = 11'd0;
wire [10:0] monroe_ionphoton_monroe_ionphoton_reader_length_storage;
reg monroe_ionphoton_monroe_ionphoton_reader_length_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_reader_irq;
wire monroe_ionphoton_monroe_ionphoton_reader_done_status;
reg monroe_ionphoton_monroe_ionphoton_reader_done_pending = 1'd0;
reg monroe_ionphoton_monroe_ionphoton_reader_done_trigger;
reg monroe_ionphoton_monroe_ionphoton_reader_done_clear;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_re;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_r;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_w;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_re;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_r;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_w;
reg monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage_full = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage;
reg monroe_ionphoton_monroe_ionphoton_reader_eventmanager_re = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_stb;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_ack;
reg monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_eop = 1'd0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_slot;
wire [10:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_length;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_source_stb;
reg monroe_ionphoton_monroe_ionphoton_reader_fifo_source_ack;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_source_eop;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_slot;
wire [10:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_we;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_re;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_readable;
wire [13:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_din;
wire [13:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_dout;
reg [2:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_level = 3'd0;
reg monroe_ionphoton_monroe_ionphoton_reader_fifo_replace = 1'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_produce = 2'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_consume = 2'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr;
wire [13:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_dat_r;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_we;
wire [13:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_dat_w;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_do_read;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_adr;
wire [13:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_dat_r;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_slot;
wire [10:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_length;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_eop;
wire [1:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_slot;
wire [10:0] monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_length;
wire monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_eop;
reg [10:0] monroe_ionphoton_monroe_ionphoton_reader_counter = 11'd0;
reg monroe_ionphoton_monroe_ionphoton_reader_counter_reset;
reg monroe_ionphoton_monroe_ionphoton_reader_counter_ce;
wire monroe_ionphoton_monroe_ionphoton_reader_last;
reg monroe_ionphoton_monroe_ionphoton_reader_last_d = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_reader_memory0_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r;
wire [8:0] monroe_ionphoton_monroe_ionphoton_reader_memory1_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r;
wire [8:0] monroe_ionphoton_monroe_ionphoton_reader_memory2_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r;
wire [8:0] monroe_ionphoton_monroe_ionphoton_reader_memory3_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r;
wire monroe_ionphoton_monroe_ionphoton_ev_irq;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_w0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_sel0;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc0;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_stb0;
reg monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_we0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_cti0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_bte0;
reg monroe_ionphoton_monroe_ionphoton_sram0_bus_err0 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram0_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_dat_r0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_w0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_sel0;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc0;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_stb0;
reg monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_we0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_cti0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_bte0;
reg monroe_ionphoton_monroe_ionphoton_sram1_bus_err0 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram1_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_dat_r0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_w0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_sel0;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc0;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_stb0;
reg monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_we0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_cti0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_bte0;
reg monroe_ionphoton_monroe_ionphoton_sram2_bus_err0 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram2_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_dat_r0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_w0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_sel0;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc0;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_stb0;
reg monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_we0;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_cti0;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_bte0;
reg monroe_ionphoton_monroe_ionphoton_sram3_bus_err0 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram3_adr0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_dat_r0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_w1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r1;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1;
reg monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram0_bus_we1;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_cti1;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram0_bus_bte1;
reg monroe_ionphoton_monroe_ionphoton_sram0_bus_err1 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram0_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_dat_r1;
reg [3:0] monroe_ionphoton_monroe_ionphoton_sram0_we;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram0_dat_w;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_w1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r1;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1;
reg monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram1_bus_we1;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_cti1;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram1_bus_bte1;
reg monroe_ionphoton_monroe_ionphoton_sram1_bus_err1 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram1_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_dat_r1;
reg [3:0] monroe_ionphoton_monroe_ionphoton_sram1_we;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram1_dat_w;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_w1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r1;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1;
reg monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram2_bus_we1;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_cti1;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram2_bus_bte1;
reg monroe_ionphoton_monroe_ionphoton_sram2_bus_err1 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram2_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_dat_r1;
reg [3:0] monroe_ionphoton_monroe_ionphoton_sram2_we;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram2_dat_w;
wire [29:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_w1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r1;
wire [3:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1;
reg monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1 = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_sram3_bus_we1;
wire [2:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_cti1;
wire [1:0] monroe_ionphoton_monroe_ionphoton_sram3_bus_bte1;
reg monroe_ionphoton_monroe_ionphoton_sram3_bus_err1 = 1'd0;
wire [8:0] monroe_ionphoton_monroe_ionphoton_sram3_adr1;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_dat_r1;
reg [3:0] monroe_ionphoton_monroe_ionphoton_sram3_we;
wire [31:0] monroe_ionphoton_monroe_ionphoton_sram3_dat_w;
reg [7:0] monroe_ionphoton_monroe_ionphoton_slave_sel;
reg [7:0] monroe_ionphoton_monroe_ionphoton_slave_sel_r = 8'd0;
reg monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage_full = 1'd1;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage;
reg monroe_ionphoton_monroe_ionphoton_kernel_cpu_re = 1'd0;
wire sys_kernel_clk;
wire sys_kernel_rst;
wire [29:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_sel;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cyc;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_stb;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_ack;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_bte;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_err;
wire [29:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_sel;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cyc;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_stb;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_ack;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_bte;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_err;
reg [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_interrupt = 32'd0;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_i_adr_o;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_d_adr_o;
wire [29:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_w;
wire [31:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_sel;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cyc;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_stb;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_ack;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_bte;
wire monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_err;
wire [29:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_sel;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i1_cyc;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i1_stb;
reg monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i1_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_mailbox_i1_bte;
reg monroe_ionphoton_monroe_ionphoton_mailbox_i1_err = 1'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_sel;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i2_cyc;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i2_stb;
reg monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_mailbox_i2_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_mailbox_i2_bte;
reg monroe_ionphoton_monroe_ionphoton_mailbox_i2_err = 1'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_mailbox0 = 32'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_mailbox1 = 32'd0;
reg [31:0] monroe_ionphoton_monroe_ionphoton_mailbox2 = 32'd0;
reg [7:0] monroe_ionphoton_add_identifier_storage_full = 8'd0;
wire [7:0] monroe_ionphoton_add_identifier_storage;
reg monroe_ionphoton_add_identifier_re = 1'd0;
wire [7:0] monroe_ionphoton_add_identifier_status;
wire [5:0] monroe_ionphoton_add_identifier_adr;
wire [7:0] monroe_ionphoton_add_identifier_dat_r;
reg monroe_ionphoton_leds_storage_full = 1'd0;
wire monroe_ionphoton_leds_storage;
reg monroe_ionphoton_leds_re = 1'd0;
reg [1:0] monroe_ionphoton_i2c_status0;
reg [1:0] monroe_ionphoton_i2c_out_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_i2c_out_storage;
reg monroe_ionphoton_i2c_out_re = 1'd0;
reg [1:0] monroe_ionphoton_i2c_oe_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_i2c_oe_storage;
reg monroe_ionphoton_i2c_oe_re = 1'd0;
wire monroe_ionphoton_i2c_tstriple0_o;
wire monroe_ionphoton_i2c_tstriple0_oe;
wire monroe_ionphoton_i2c_tstriple0_i;
wire monroe_ionphoton_i2c_status1;
wire monroe_ionphoton_i2c_tstriple1_o;
wire monroe_ionphoton_i2c_tstriple1_oe;
wire monroe_ionphoton_i2c_tstriple1_i;
wire monroe_ionphoton_i2c_status2;
reg [7:0] inout_8x0_serdes_o0 = 8'd0;
wire [7:0] inout_8x0_serdes_i0;
reg inout_8x0_serdes_oe = 1'd0;
wire inout_8x0_serdes_pad_i0;
wire inout_8x0_serdes_pad_o0;
wire [7:0] inout_8x0_serdes_i1;
wire inout_8x0_serdes_pad_i1;
wire [7:0] inout_8x0_serdes_o1;
wire inout_8x0_serdes_t_in;
wire inout_8x0_serdes_t_out;
wire inout_8x0_serdes_pad_o1;
reg inout_8x0_inout_8x0_ointerface0_stb = 1'd0;
reg inout_8x0_inout_8x0_ointerface0_busy = 1'd0;
reg [1:0] inout_8x0_inout_8x0_ointerface0_data = 2'd0;
reg [1:0] inout_8x0_inout_8x0_ointerface0_address = 2'd0;
reg [2:0] inout_8x0_inout_8x0_ointerface0_fine_ts = 3'd0;
reg inout_8x0_inout_8x0_iinterface0_stb = 1'd0;
reg inout_8x0_inout_8x0_iinterface0_data = 1'd0;
reg [2:0] inout_8x0_inout_8x0_iinterface0_fine_ts = 3'd0;
wire inout_8x0_inout_8x0_override_en;
wire inout_8x0_inout_8x0_override_o;
wire inout_8x0_inout_8x0_override_oe;
wire inout_8x0_inout_8x0_input_state;
reg inout_8x0_inout_8x0_previous_data = 1'd0;
reg inout_8x0_inout_8x0_oe_k = 1'd0;
reg [1:0] inout_8x0_inout_8x0_sensitivity = 2'd0;
reg inout_8x0_inout_8x0_sample = 1'd0;
reg inout_8x0_inout_8x0_i_d = 1'd0;
wire [7:0] inout_8x0_inout_8x0_i;
reg [2:0] inout_8x0_inout_8x0_o;
wire inout_8x0_inout_8x0_n;
reg [7:0] inout_8x1_serdes_o0 = 8'd0;
wire [7:0] inout_8x1_serdes_i0;
reg inout_8x1_serdes_oe = 1'd0;
wire inout_8x1_serdes_pad_i0;
wire inout_8x1_serdes_pad_o0;
wire [7:0] inout_8x1_serdes_i1;
wire inout_8x1_serdes_pad_i1;
wire [7:0] inout_8x1_serdes_o1;
wire inout_8x1_serdes_t_in;
wire inout_8x1_serdes_t_out;
wire inout_8x1_serdes_pad_o1;
reg inout_8x1_inout_8x1_ointerface1_stb = 1'd0;
reg inout_8x1_inout_8x1_ointerface1_busy = 1'd0;
reg [1:0] inout_8x1_inout_8x1_ointerface1_data = 2'd0;
reg [1:0] inout_8x1_inout_8x1_ointerface1_address = 2'd0;
reg [2:0] inout_8x1_inout_8x1_ointerface1_fine_ts = 3'd0;
reg inout_8x1_inout_8x1_iinterface1_stb = 1'd0;
reg inout_8x1_inout_8x1_iinterface1_data = 1'd0;
reg [2:0] inout_8x1_inout_8x1_iinterface1_fine_ts = 3'd0;
wire inout_8x1_inout_8x1_override_en;
wire inout_8x1_inout_8x1_override_o;
wire inout_8x1_inout_8x1_override_oe;
wire inout_8x1_inout_8x1_input_state;
reg inout_8x1_inout_8x1_previous_data = 1'd0;
reg inout_8x1_inout_8x1_oe_k = 1'd0;
reg [1:0] inout_8x1_inout_8x1_sensitivity = 2'd0;
reg inout_8x1_inout_8x1_sample = 1'd0;
reg inout_8x1_inout_8x1_i_d = 1'd0;
wire [7:0] inout_8x1_inout_8x1_i;
reg [2:0] inout_8x1_inout_8x1_o;
wire inout_8x1_inout_8x1_n;
reg [7:0] inout_8x2_serdes_o0 = 8'd0;
wire [7:0] inout_8x2_serdes_i0;
reg inout_8x2_serdes_oe = 1'd0;
wire inout_8x2_serdes_pad_i0;
wire inout_8x2_serdes_pad_o0;
wire [7:0] inout_8x2_serdes_i1;
wire inout_8x2_serdes_pad_i1;
wire [7:0] inout_8x2_serdes_o1;
wire inout_8x2_serdes_t_in;
wire inout_8x2_serdes_t_out;
wire inout_8x2_serdes_pad_o1;
reg inout_8x2_inout_8x2_ointerface2_stb = 1'd0;
reg inout_8x2_inout_8x2_ointerface2_busy = 1'd0;
reg [1:0] inout_8x2_inout_8x2_ointerface2_data = 2'd0;
reg [1:0] inout_8x2_inout_8x2_ointerface2_address = 2'd0;
reg [2:0] inout_8x2_inout_8x2_ointerface2_fine_ts = 3'd0;
reg inout_8x2_inout_8x2_iinterface2_stb = 1'd0;
reg inout_8x2_inout_8x2_iinterface2_data = 1'd0;
reg [2:0] inout_8x2_inout_8x2_iinterface2_fine_ts = 3'd0;
wire inout_8x2_inout_8x2_override_en;
wire inout_8x2_inout_8x2_override_o;
wire inout_8x2_inout_8x2_override_oe;
wire inout_8x2_inout_8x2_input_state;
reg inout_8x2_inout_8x2_previous_data = 1'd0;
reg inout_8x2_inout_8x2_oe_k = 1'd0;
reg [1:0] inout_8x2_inout_8x2_sensitivity = 2'd0;
reg inout_8x2_inout_8x2_sample = 1'd0;
reg inout_8x2_inout_8x2_i_d = 1'd0;
wire [7:0] inout_8x2_inout_8x2_i;
reg [2:0] inout_8x2_inout_8x2_o;
wire inout_8x2_inout_8x2_n;
reg [7:0] inout_8x3_serdes_o0 = 8'd0;
wire [7:0] inout_8x3_serdes_i0;
reg inout_8x3_serdes_oe = 1'd0;
wire inout_8x3_serdes_pad_i0;
wire inout_8x3_serdes_pad_o0;
wire [7:0] inout_8x3_serdes_i1;
wire inout_8x3_serdes_pad_i1;
wire [7:0] inout_8x3_serdes_o1;
wire inout_8x3_serdes_t_in;
wire inout_8x3_serdes_t_out;
wire inout_8x3_serdes_pad_o1;
reg inout_8x3_inout_8x3_ointerface3_stb = 1'd0;
reg inout_8x3_inout_8x3_ointerface3_busy = 1'd0;
reg [1:0] inout_8x3_inout_8x3_ointerface3_data = 2'd0;
reg [1:0] inout_8x3_inout_8x3_ointerface3_address = 2'd0;
reg [2:0] inout_8x3_inout_8x3_ointerface3_fine_ts = 3'd0;
reg inout_8x3_inout_8x3_iinterface3_stb = 1'd0;
reg inout_8x3_inout_8x3_iinterface3_data = 1'd0;
reg [2:0] inout_8x3_inout_8x3_iinterface3_fine_ts = 3'd0;
wire inout_8x3_inout_8x3_override_en;
wire inout_8x3_inout_8x3_override_o;
wire inout_8x3_inout_8x3_override_oe;
wire inout_8x3_inout_8x3_input_state;
reg inout_8x3_inout_8x3_previous_data = 1'd0;
reg inout_8x3_inout_8x3_oe_k = 1'd0;
reg [1:0] inout_8x3_inout_8x3_sensitivity = 2'd0;
reg inout_8x3_inout_8x3_sample = 1'd0;
reg inout_8x3_inout_8x3_i_d = 1'd0;
wire [7:0] inout_8x3_inout_8x3_i;
reg [2:0] inout_8x3_inout_8x3_o;
wire inout_8x3_inout_8x3_n;
reg [7:0] output_8x0_o = 8'd0;
reg output_8x0_t_in = 1'd0;
wire output_8x0_t_out;
wire output_8x0_pad_o;
reg output_8x0_stb = 1'd0;
reg output_8x0_busy = 1'd0;
reg output_8x0_data = 1'd0;
reg [2:0] output_8x0_fine_ts = 3'd0;
wire output_8x0_override_en;
wire output_8x0_override_o;
reg output_8x0_previous_data = 1'd0;
reg [7:0] output_8x1_o = 8'd0;
reg output_8x1_t_in = 1'd0;
wire output_8x1_t_out;
wire output_8x1_pad_o;
reg output_8x1_stb = 1'd0;
reg output_8x1_busy = 1'd0;
reg output_8x1_data = 1'd0;
reg [2:0] output_8x1_fine_ts = 3'd0;
wire output_8x1_override_en;
wire output_8x1_override_o;
reg output_8x1_previous_data = 1'd0;
reg [7:0] output_8x2_o = 8'd0;
reg output_8x2_t_in = 1'd0;
wire output_8x2_t_out;
wire output_8x2_pad_o;
reg output_8x2_stb = 1'd0;
reg output_8x2_busy = 1'd0;
reg output_8x2_data = 1'd0;
reg [2:0] output_8x2_fine_ts = 3'd0;
wire output_8x2_override_en;
wire output_8x2_override_o;
reg output_8x2_previous_data = 1'd0;
reg [7:0] output_8x3_o = 8'd0;
reg output_8x3_t_in = 1'd0;
wire output_8x3_t_out;
wire output_8x3_pad_o;
reg output_8x3_stb = 1'd0;
reg output_8x3_busy = 1'd0;
reg output_8x3_data = 1'd0;
reg [2:0] output_8x3_fine_ts = 3'd0;
wire output_8x3_override_en;
wire output_8x3_override_o;
reg output_8x3_previous_data = 1'd0;
reg [7:0] output_8x4_o = 8'd0;
reg output_8x4_t_in = 1'd0;
wire output_8x4_t_out;
wire output_8x4_pad_o;
reg output_8x4_stb = 1'd0;
reg output_8x4_busy = 1'd0;
reg output_8x4_data = 1'd0;
reg [2:0] output_8x4_fine_ts = 3'd0;
wire output_8x4_override_en;
wire output_8x4_override_o;
reg output_8x4_previous_data = 1'd0;
reg [7:0] output_8x5_o = 8'd0;
reg output_8x5_t_in = 1'd0;
wire output_8x5_t_out;
wire output_8x5_pad_o;
reg output_8x5_stb = 1'd0;
reg output_8x5_busy = 1'd0;
reg output_8x5_data = 1'd0;
reg [2:0] output_8x5_fine_ts = 3'd0;
wire output_8x5_override_en;
wire output_8x5_override_o;
reg output_8x5_previous_data = 1'd0;
reg [7:0] output_8x6_o = 8'd0;
reg output_8x6_t_in = 1'd0;
wire output_8x6_t_out;
wire output_8x6_pad_o;
reg output_8x6_stb = 1'd0;
reg output_8x6_busy = 1'd0;
reg output_8x6_data = 1'd0;
reg [2:0] output_8x6_fine_ts = 3'd0;
wire output_8x6_override_en;
wire output_8x6_override_o;
reg output_8x6_previous_data = 1'd0;
reg [7:0] output_8x7_o = 8'd0;
reg output_8x7_t_in = 1'd0;
wire output_8x7_t_out;
wire output_8x7_pad_o;
reg output_8x7_stb = 1'd0;
reg output_8x7_busy = 1'd0;
reg output_8x7_data = 1'd0;
reg [2:0] output_8x7_fine_ts = 3'd0;
wire output_8x7_override_en;
wire output_8x7_override_o;
reg output_8x7_previous_data = 1'd0;
reg [7:0] output_8x8_o = 8'd0;
reg output_8x8_t_in = 1'd0;
wire output_8x8_t_out;
wire output_8x8_pad_o;
reg output_8x8_stb = 1'd0;
reg output_8x8_busy = 1'd0;
reg output_8x8_data = 1'd0;
reg [2:0] output_8x8_fine_ts = 3'd0;
wire output_8x8_override_en;
wire output_8x8_override_o;
reg output_8x8_previous_data = 1'd0;
reg [7:0] output_8x9_o = 8'd0;
reg output_8x9_t_in = 1'd0;
wire output_8x9_t_out;
wire output_8x9_pad_o;
reg output_8x9_stb = 1'd0;
reg output_8x9_busy = 1'd0;
reg output_8x9_data = 1'd0;
reg [2:0] output_8x9_fine_ts = 3'd0;
wire output_8x9_override_en;
wire output_8x9_override_o;
reg output_8x9_previous_data = 1'd0;
reg [7:0] output_8x10_o = 8'd0;
reg output_8x10_t_in = 1'd0;
wire output_8x10_t_out;
wire output_8x10_pad_o;
reg output_8x10_stb = 1'd0;
reg output_8x10_busy = 1'd0;
reg output_8x10_data = 1'd0;
reg [2:0] output_8x10_fine_ts = 3'd0;
wire output_8x10_override_en;
wire output_8x10_override_o;
reg output_8x10_previous_data = 1'd0;
reg [7:0] output_8x11_o = 8'd0;
reg output_8x11_t_in = 1'd0;
wire output_8x11_t_out;
wire output_8x11_pad_o;
reg output_8x11_stb = 1'd0;
reg output_8x11_busy = 1'd0;
reg output_8x11_data = 1'd0;
reg [2:0] output_8x11_fine_ts = 3'd0;
wire output_8x11_override_en;
wire output_8x11_override_o;
reg output_8x11_previous_data = 1'd0;
wire [2:0] spimaster0_interface_cs0;
wire [2:0] spimaster0_interface_cs_polarity;
wire spimaster0_interface_clk_next;
wire spimaster0_interface_clk_polarity;
wire spimaster0_interface_cs_next;
wire spimaster0_interface_ce;
wire spimaster0_interface_sample;
wire spimaster0_interface_offline;
wire spimaster0_interface_half_duplex;
wire spimaster0_interface_sdi;
wire spimaster0_interface_sdo;
reg [2:0] spimaster0_interface_cs1 = 3'd7;
reg spimaster0_interface_clk = 1'd0;
wire spimaster0_interface_miso;
wire spimaster0_interface_mosi;
reg spimaster0_interface_miso_reg = 1'd0;
reg spimaster0_interface_mosi_reg = 1'd0;
wire [4:0] spimaster0_spimachine0_length;
wire spimaster0_spimachine0_clk_phase;
reg spimaster0_spimachine0_clk_next;
reg spimaster0_spimachine0_cs_next;
wire spimaster0_spimachine0_ce;
reg spimaster0_spimachine0_idle;
wire spimaster0_spimachine0_load0;
reg spimaster0_spimachine0_readable;
reg spimaster0_spimachine0_writable;
wire spimaster0_spimachine0_end0;
wire [31:0] spimaster0_spimachine0_pdo;
wire [31:0] spimaster0_spimachine0_pdi;
reg spimaster0_spimachine0_sdo = 1'd0;
wire spimaster0_spimachine0_sdi;
wire spimaster0_spimachine0_lsb_first;
reg spimaster0_spimachine0_load1;
reg spimaster0_spimachine0_shift;
reg spimaster0_spimachine0_sample;
reg [31:0] spimaster0_spimachine0_sr = 32'd0;
wire [7:0] spimaster0_spimachine0_div;
reg spimaster0_spimachine0_extend;
wire spimaster0_spimachine0_done;
reg spimaster0_spimachine0_count;
reg [6:0] spimaster0_spimachine0_cnt = 7'd0;
wire spimaster0_spimachine0_cnt_done;
reg spimaster0_spimachine0_do_extend = 1'd0;
reg [4:0] spimaster0_spimachine0_n = 5'd0;
reg spimaster0_spimachine0_end1 = 1'd0;
reg spimaster0_ointerface0_stb = 1'd0;
wire spimaster0_ointerface0_busy;
reg [31:0] spimaster0_ointerface0_data = 32'd0;
reg spimaster0_ointerface0_address = 1'd0;
wire spimaster0_iinterface0_stb;
wire [31:0] spimaster0_iinterface0_data;
reg spimaster0_config_offline = 1'd1;
reg spimaster0_config_end = 1'd1;
reg spimaster0_config_input = 1'd0;
reg spimaster0_config_cs_polarity = 1'd0;
reg spimaster0_config_clk_polarity = 1'd0;
reg spimaster0_config_clk_phase = 1'd0;
reg spimaster0_config_lsb_first = 1'd0;
reg spimaster0_config_half_duplex = 1'd0;
reg [4:0] spimaster0_config_length = 5'd0;
reg [2:0] spimaster0_config_padding = 3'd0;
reg [7:0] spimaster0_config_div = 8'd0;
reg [7:0] spimaster0_config_cs = 8'd0;
reg spimaster0_read = 1'd0;
reg pad0 = 1'd0;
reg [7:0] output_8x12_o = 8'd0;
reg output_8x12_t_in = 1'd0;
wire output_8x12_t_out;
wire output_8x12_pad_o;
reg output_8x12_stb = 1'd0;
reg output_8x12_busy = 1'd0;
reg output_8x12_data = 1'd0;
reg [2:0] output_8x12_fine_ts = 3'd0;
wire output_8x12_override_en;
wire output_8x12_override_o;
reg output_8x12_previous_data = 1'd0;
reg [7:0] output_8x13_o = 8'd0;
reg output_8x13_t_in = 1'd0;
wire output_8x13_t_out;
wire output_8x13_pad_o;
reg output_8x13_stb = 1'd0;
reg output_8x13_busy = 1'd0;
reg output_8x13_data = 1'd0;
reg [2:0] output_8x13_fine_ts = 3'd0;
wire output_8x13_override_en;
wire output_8x13_override_o;
reg output_8x13_previous_data = 1'd0;
reg [7:0] output_8x14_o = 8'd0;
reg output_8x14_t_in = 1'd0;
wire output_8x14_t_out;
wire output_8x14_pad_o;
reg output_8x14_stb = 1'd0;
reg output_8x14_busy = 1'd0;
reg output_8x14_data = 1'd0;
reg [2:0] output_8x14_fine_ts = 3'd0;
wire output_8x14_override_en;
wire output_8x14_override_o;
reg output_8x14_previous_data = 1'd0;
reg [7:0] output_8x15_o = 8'd0;
reg output_8x15_t_in = 1'd0;
wire output_8x15_t_out;
wire output_8x15_pad_o;
reg output_8x15_stb = 1'd0;
reg output_8x15_busy = 1'd0;
reg output_8x15_data = 1'd0;
reg [2:0] output_8x15_fine_ts = 3'd0;
wire output_8x15_override_en;
wire output_8x15_override_o;
reg output_8x15_previous_data = 1'd0;
reg [7:0] output_8x16_o = 8'd0;
reg output_8x16_t_in = 1'd0;
wire output_8x16_t_out;
wire output_8x16_pad_o;
reg output_8x16_stb = 1'd0;
reg output_8x16_busy = 1'd0;
reg output_8x16_data = 1'd0;
reg [2:0] output_8x16_fine_ts = 3'd0;
wire output_8x16_override_en;
wire output_8x16_override_o;
reg output_8x16_previous_data = 1'd0;
wire [2:0] spimaster1_interface_cs0;
wire [2:0] spimaster1_interface_cs_polarity;
wire spimaster1_interface_clk_next;
wire spimaster1_interface_clk_polarity;
wire spimaster1_interface_cs_next;
wire spimaster1_interface_ce;
wire spimaster1_interface_sample;
wire spimaster1_interface_offline;
wire spimaster1_interface_half_duplex;
wire spimaster1_interface_sdi;
wire spimaster1_interface_sdo;
reg [2:0] spimaster1_interface_cs1 = 3'd7;
reg spimaster1_interface_clk = 1'd0;
wire spimaster1_interface_miso;
wire spimaster1_interface_mosi;
reg spimaster1_interface_miso_reg = 1'd0;
reg spimaster1_interface_mosi_reg = 1'd0;
wire [4:0] spimaster1_spimachine1_length;
wire spimaster1_spimachine1_clk_phase;
reg spimaster1_spimachine1_clk_next;
reg spimaster1_spimachine1_cs_next;
wire spimaster1_spimachine1_ce;
reg spimaster1_spimachine1_idle;
wire spimaster1_spimachine1_load0;
reg spimaster1_spimachine1_readable;
reg spimaster1_spimachine1_writable;
wire spimaster1_spimachine1_end0;
wire [31:0] spimaster1_spimachine1_pdo;
wire [31:0] spimaster1_spimachine1_pdi;
reg spimaster1_spimachine1_sdo = 1'd0;
wire spimaster1_spimachine1_sdi;
wire spimaster1_spimachine1_lsb_first;
reg spimaster1_spimachine1_load1;
reg spimaster1_spimachine1_shift;
reg spimaster1_spimachine1_sample;
reg [31:0] spimaster1_spimachine1_sr = 32'd0;
wire [7:0] spimaster1_spimachine1_div;
reg spimaster1_spimachine1_extend;
wire spimaster1_spimachine1_done;
reg spimaster1_spimachine1_count;
reg [6:0] spimaster1_spimachine1_cnt = 7'd0;
wire spimaster1_spimachine1_cnt_done;
reg spimaster1_spimachine1_do_extend = 1'd0;
reg [4:0] spimaster1_spimachine1_n = 5'd0;
reg spimaster1_spimachine1_end1 = 1'd0;
reg spimaster1_ointerface1_stb = 1'd0;
wire spimaster1_ointerface1_busy;
reg [31:0] spimaster1_ointerface1_data = 32'd0;
reg spimaster1_ointerface1_address = 1'd0;
wire spimaster1_iinterface1_stb;
wire [31:0] spimaster1_iinterface1_data;
reg spimaster1_config_offline = 1'd1;
reg spimaster1_config_end = 1'd1;
reg spimaster1_config_input = 1'd0;
reg spimaster1_config_cs_polarity = 1'd0;
reg spimaster1_config_clk_polarity = 1'd0;
reg spimaster1_config_clk_phase = 1'd0;
reg spimaster1_config_lsb_first = 1'd0;
reg spimaster1_config_half_duplex = 1'd0;
reg [4:0] spimaster1_config_length = 5'd0;
reg [2:0] spimaster1_config_padding = 3'd0;
reg [7:0] spimaster1_config_div = 8'd0;
reg [7:0] spimaster1_config_cs = 8'd0;
reg spimaster1_read = 1'd0;
reg pad1 = 1'd0;
reg [7:0] output_8x17_o = 8'd0;
reg output_8x17_t_in = 1'd0;
wire output_8x17_t_out;
wire output_8x17_pad_o;
reg output_8x17_stb = 1'd0;
reg output_8x17_busy = 1'd0;
reg output_8x17_data = 1'd0;
reg [2:0] output_8x17_fine_ts = 3'd0;
wire output_8x17_override_en;
wire output_8x17_override_o;
reg output_8x17_previous_data = 1'd0;
reg [7:0] output_8x18_o = 8'd0;
reg output_8x18_t_in = 1'd0;
wire output_8x18_t_out;
wire output_8x18_pad_o;
reg output_8x18_stb = 1'd0;
reg output_8x18_busy = 1'd0;
reg output_8x18_data = 1'd0;
reg [2:0] output_8x18_fine_ts = 3'd0;
wire output_8x18_override_en;
wire output_8x18_override_o;
reg output_8x18_previous_data = 1'd0;
reg [7:0] output_8x19_o = 8'd0;
reg output_8x19_t_in = 1'd0;
wire output_8x19_t_out;
wire output_8x19_pad_o;
reg output_8x19_stb = 1'd0;
reg output_8x19_busy = 1'd0;
reg output_8x19_data = 1'd0;
reg [2:0] output_8x19_fine_ts = 3'd0;
wire output_8x19_override_en;
wire output_8x19_override_o;
reg output_8x19_previous_data = 1'd0;
reg [7:0] output_8x20_o = 8'd0;
reg output_8x20_t_in = 1'd0;
wire output_8x20_t_out;
wire output_8x20_pad_o;
reg output_8x20_stb = 1'd0;
reg output_8x20_busy = 1'd0;
reg output_8x20_data = 1'd0;
reg [2:0] output_8x20_fine_ts = 3'd0;
wire output_8x20_override_en;
wire output_8x20_override_o;
reg output_8x20_previous_data = 1'd0;
reg [7:0] output_8x21_o = 8'd0;
reg output_8x21_t_in = 1'd0;
wire output_8x21_t_out;
wire output_8x21_pad_o;
reg output_8x21_stb = 1'd0;
reg output_8x21_busy = 1'd0;
reg output_8x21_data = 1'd0;
reg [2:0] output_8x21_fine_ts = 3'd0;
wire output_8x21_override_en;
wire output_8x21_override_o;
reg output_8x21_previous_data = 1'd0;
wire [2:0] spimaster2_interface_cs0;
wire [2:0] spimaster2_interface_cs_polarity;
wire spimaster2_interface_clk_next;
wire spimaster2_interface_clk_polarity;
wire spimaster2_interface_cs_next;
wire spimaster2_interface_ce;
wire spimaster2_interface_sample;
wire spimaster2_interface_offline;
wire spimaster2_interface_half_duplex;
wire spimaster2_interface_sdi;
wire spimaster2_interface_sdo;
reg [2:0] spimaster2_interface_cs1 = 3'd7;
reg spimaster2_interface_clk = 1'd0;
wire spimaster2_interface_miso;
wire spimaster2_interface_mosi;
reg spimaster2_interface_miso_reg = 1'd0;
reg spimaster2_interface_mosi_reg = 1'd0;
wire [4:0] spimaster2_spimachine2_length;
wire spimaster2_spimachine2_clk_phase;
reg spimaster2_spimachine2_clk_next;
reg spimaster2_spimachine2_cs_next;
wire spimaster2_spimachine2_ce;
reg spimaster2_spimachine2_idle;
wire spimaster2_spimachine2_load0;
reg spimaster2_spimachine2_readable;
reg spimaster2_spimachine2_writable;
wire spimaster2_spimachine2_end0;
wire [31:0] spimaster2_spimachine2_pdo;
wire [31:0] spimaster2_spimachine2_pdi;
reg spimaster2_spimachine2_sdo = 1'd0;
wire spimaster2_spimachine2_sdi;
wire spimaster2_spimachine2_lsb_first;
reg spimaster2_spimachine2_load1;
reg spimaster2_spimachine2_shift;
reg spimaster2_spimachine2_sample;
reg [31:0] spimaster2_spimachine2_sr = 32'd0;
wire [7:0] spimaster2_spimachine2_div;
reg spimaster2_spimachine2_extend;
wire spimaster2_spimachine2_done;
reg spimaster2_spimachine2_count;
reg [6:0] spimaster2_spimachine2_cnt = 7'd0;
wire spimaster2_spimachine2_cnt_done;
reg spimaster2_spimachine2_do_extend = 1'd0;
reg [4:0] spimaster2_spimachine2_n = 5'd0;
reg spimaster2_spimachine2_end1 = 1'd0;
reg spimaster2_ointerface2_stb = 1'd0;
wire spimaster2_ointerface2_busy;
reg [31:0] spimaster2_ointerface2_data = 32'd0;
reg spimaster2_ointerface2_address = 1'd0;
wire spimaster2_iinterface2_stb;
wire [31:0] spimaster2_iinterface2_data;
reg spimaster2_config_offline = 1'd1;
reg spimaster2_config_end = 1'd1;
reg spimaster2_config_input = 1'd0;
reg spimaster2_config_cs_polarity = 1'd0;
reg spimaster2_config_clk_polarity = 1'd0;
reg spimaster2_config_clk_phase = 1'd0;
reg spimaster2_config_lsb_first = 1'd0;
reg spimaster2_config_half_duplex = 1'd0;
reg [4:0] spimaster2_config_length = 5'd0;
reg [2:0] spimaster2_config_padding = 3'd0;
reg [7:0] spimaster2_config_div = 8'd0;
reg [7:0] spimaster2_config_cs = 8'd0;
reg spimaster2_read = 1'd0;
reg pad2 = 1'd0;
reg [7:0] output_8x22_o = 8'd0;
reg output_8x22_t_in = 1'd0;
wire output_8x22_t_out;
wire output_8x22_pad_o;
reg output_8x22_stb = 1'd0;
reg output_8x22_busy = 1'd0;
reg output_8x22_data = 1'd0;
reg [2:0] output_8x22_fine_ts = 3'd0;
wire output_8x22_override_en;
wire output_8x22_override_o;
reg output_8x22_previous_data = 1'd0;
reg [7:0] output_8x23_o = 8'd0;
reg output_8x23_t_in = 1'd0;
wire output_8x23_t_out;
wire output_8x23_pad_o;
reg output_8x23_stb = 1'd0;
reg output_8x23_busy = 1'd0;
reg output_8x23_data = 1'd0;
reg [2:0] output_8x23_fine_ts = 3'd0;
wire output_8x23_override_en;
wire output_8x23_override_o;
reg output_8x23_previous_data = 1'd0;
reg [7:0] output_8x24_o = 8'd0;
reg output_8x24_t_in = 1'd0;
wire output_8x24_t_out;
wire output_8x24_pad_o;
reg output_8x24_stb = 1'd0;
reg output_8x24_busy = 1'd0;
reg output_8x24_data = 1'd0;
reg [2:0] output_8x24_fine_ts = 3'd0;
wire output_8x24_override_en;
wire output_8x24_override_o;
reg output_8x24_previous_data = 1'd0;
reg [7:0] output_8x25_o = 8'd0;
reg output_8x25_t_in = 1'd0;
wire output_8x25_t_out;
wire output_8x25_pad_o;
reg output_8x25_stb = 1'd0;
reg output_8x25_busy = 1'd0;
reg output_8x25_data = 1'd0;
reg [2:0] output_8x25_fine_ts = 3'd0;
wire output_8x25_override_en;
wire output_8x25_override_o;
reg output_8x25_previous_data = 1'd0;
reg [7:0] output_8x26_o = 8'd0;
reg output_8x26_t_in = 1'd0;
wire output_8x26_t_out;
wire output_8x26_pad_o;
reg output_8x26_stb = 1'd0;
reg output_8x26_busy = 1'd0;
reg output_8x26_data = 1'd0;
reg [2:0] output_8x26_fine_ts = 3'd0;
wire output_8x26_override_en;
wire output_8x26_override_o;
reg output_8x26_previous_data = 1'd0;
reg output0_stb = 1'd0;
reg output0_busy = 1'd0;
reg output0_data = 1'd0;
reg output0_pad_o = 1'd0;
wire output0_override_en;
wire output0_override_o;
reg output0_pad_k = 1'd0;
reg output1_stb = 1'd0;
reg output1_busy = 1'd0;
reg output1_data = 1'd0;
reg output1_pad_o = 1'd0;
wire output1_override_en;
wire output1_override_o;
reg output1_pad_k = 1'd0;
reg stb = 1'd0;
reg busy = 1'd0;
reg [31:0] data = 32'd0;
reg monroe_ionphoton_rtio_crg_storage_full = 1'd1;
wire monroe_ionphoton_rtio_crg_storage;
reg monroe_ionphoton_rtio_crg_re = 1'd0;
wire monroe_ionphoton_rtio_crg_pll_locked_status;
wire rtio_clk;
wire rtio_rst;
wire rtiox4_clk;
wire monroe_ionphoton_rtio_crg_clk_synth_se;
wire monroe_ionphoton_rtio_crg_pll_locked;
wire monroe_ionphoton_rtio_crg_rtio_clk;
wire monroe_ionphoton_rtio_crg_rtiox4_clk;
wire monroe_ionphoton_rtio_crg_fb_clk;
reg [60:0] monroe_ionphoton_rtio_tsc_coarse_ts = 61'd0;
wire [63:0] monroe_ionphoton_rtio_tsc_full_ts;
wire [60:0] monroe_ionphoton_rtio_tsc_coarse_ts_sys;
wire [63:0] monroe_ionphoton_rtio_tsc_full_ts_sys;
reg monroe_ionphoton_rtio_tsc_load = 1'd0;
reg [60:0] monroe_ionphoton_rtio_tsc_load_value = 61'd0;
wire [60:0] monroe_ionphoton_rtio_tsc_i;
reg [60:0] monroe_ionphoton_rtio_tsc_o = 61'd0;
(* dont_touch = "true" *) reg [60:0] monroe_ionphoton_rtio_tsc_value_gray_rtio = 61'd0;
wire [60:0] monroe_ionphoton_rtio_tsc_value_gray_sys;
reg [60:0] monroe_ionphoton_rtio_tsc_value_sys;
reg [1:0] monroe_ionphoton_rtio_core_cri_cmd;
wire [23:0] monroe_ionphoton_rtio_core_cri_chan_sel;
wire [63:0] monroe_ionphoton_rtio_core_cri_o_timestamp;
wire [511:0] monroe_ionphoton_rtio_core_cri_o_data;
wire [7:0] monroe_ionphoton_rtio_core_cri_o_address;
wire [2:0] monroe_ionphoton_rtio_core_cri_o_status;
reg monroe_ionphoton_rtio_core_cri_o_buffer_space_valid = 1'd0;
reg [15:0] monroe_ionphoton_rtio_core_cri_o_buffer_space = 16'd0;
wire [63:0] monroe_ionphoton_rtio_core_cri_i_timeout;
reg [31:0] monroe_ionphoton_rtio_core_cri_i_data = 32'd0;
reg [63:0] monroe_ionphoton_rtio_core_cri_i_timestamp = 64'd0;
reg [3:0] monroe_ionphoton_rtio_core_cri_i_status = 4'd0;
wire monroe_ionphoton_rtio_core_reset_re;
wire monroe_ionphoton_rtio_core_reset_r;
reg monroe_ionphoton_rtio_core_reset_w = 1'd0;
wire monroe_ionphoton_rtio_core_reset_phy_re;
wire monroe_ionphoton_rtio_core_reset_phy_r;
reg monroe_ionphoton_rtio_core_reset_phy_w = 1'd0;
wire monroe_ionphoton_rtio_core_async_error_re;
wire [2:0] monroe_ionphoton_rtio_core_async_error_r;
wire [2:0] monroe_ionphoton_rtio_core_async_error_w;
reg [15:0] monroe_ionphoton_rtio_core_collision_channel_status = 16'd0;
reg [15:0] monroe_ionphoton_rtio_core_busy_channel_status = 16'd0;
reg [15:0] monroe_ionphoton_rtio_core_sequence_error_channel_status = 16'd0;
(* dont_touch = "true" *) reg monroe_ionphoton_rtio_core_cmd_reset = 1'd1;
(* dont_touch = "true" *) reg monroe_ionphoton_rtio_core_cmd_reset_phy = 1'd1;
wire rsys_clk;
wire rsys_rst;
wire rio_clk;
wire rio_rst;
wire rio_phy_clk;
wire rio_phy_rst;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error = 1'd0;
reg [15:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error_channel = 16'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp = 61'd0;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_data;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_we;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_seqn;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_channel;
reg [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_address;
wire [31:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_data;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_wait;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_underflow = 1'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane = 3'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_coarse_timestamp = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 = 61'd0;
reg [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 = 61'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn = 12'd0;
wire [60:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp;
reg signed [61:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_min_minus_timestamp = 62'sd0;
reg signed [61:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp = 62'sd0;
reg signed [61:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp = 62'sd0;
reg signed [61:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_last_minus_timestamp = 62'sd0;
wire [2:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_plus_one;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_quash = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_adr;
wire [13:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_dat_r;
wire signed [13:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_min;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_last;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_lane_min;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_force_laneB = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_use_laneB;
reg [2:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_do_underflow;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_do_sequence_error;
wire [63:0] monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
wire monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable;
reg monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable_r = 1'd1;
wire monroe_ionphoton_rtio_core_outputs_record0_we;
wire monroe_ionphoton_rtio_core_outputs_record0_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record0_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record0_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record0_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record0_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record1_we;
wire monroe_ionphoton_rtio_core_outputs_record1_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record1_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record1_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record1_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record1_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record2_we;
wire monroe_ionphoton_rtio_core_outputs_record2_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record2_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record2_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record2_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record2_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record3_we;
wire monroe_ionphoton_rtio_core_outputs_record3_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record3_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record3_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record3_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record3_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record4_we;
wire monroe_ionphoton_rtio_core_outputs_record4_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record4_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record4_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record4_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record4_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record5_we;
wire monroe_ionphoton_rtio_core_outputs_record5_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record5_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record5_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record5_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record5_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record6_we;
wire monroe_ionphoton_rtio_core_outputs_record6_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record6_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record6_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record6_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record6_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record7_we;
wire monroe_ionphoton_rtio_core_outputs_record7_writable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record7_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record7_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record7_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record7_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_record0_re;
wire monroe_ionphoton_rtio_core_outputs_record0_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record0_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record0_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record0_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record0_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record1_re;
wire monroe_ionphoton_rtio_core_outputs_record1_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record1_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record1_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record1_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record1_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record2_re;
wire monroe_ionphoton_rtio_core_outputs_record2_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record2_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record2_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record2_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record2_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record3_re;
wire monroe_ionphoton_rtio_core_outputs_record3_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record3_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record3_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record3_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record3_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record4_re;
wire monroe_ionphoton_rtio_core_outputs_record4_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record4_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record4_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record4_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record4_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record5_re;
wire monroe_ionphoton_rtio_core_outputs_record5_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record5_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record5_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record5_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record5_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record6_re;
wire monroe_ionphoton_rtio_core_outputs_record6_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record6_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record6_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record6_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record6_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_record7_re;
wire monroe_ionphoton_rtio_core_outputs_record7_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record7_seqn1;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record7_payload_channel1;
wire [63:0] monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp1;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record7_payload_address1;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record7_payload_data1;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_re;
reg monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable = 1'd0;
reg [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_dout = 116'd0;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce;
(* dont_touch = "true" *) reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q = 8'd0;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary = 8'd0;
reg [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_produce_rdomain;
wire [7:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_consume_wdomain;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_we;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
wire [6:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
wire [115:0] monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;
wire monroe_ionphoton_rtio_core_outputs_gates_record0_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record0_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record0_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record1_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record1_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record1_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record2_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record2_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record2_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record3_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record3_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record3_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record4_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record4_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record4_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record5_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record5_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record5_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record6_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record6_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record6_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data0;
wire monroe_ionphoton_rtio_core_outputs_gates_record7_re;
wire monroe_ionphoton_rtio_core_outputs_gates_record7_readable;
wire [11:0] monroe_ionphoton_rtio_core_outputs_gates_record7_seqn0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel0;
wire [63:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_timestamp;
wire [1:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address0;
wire [31:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data0;
reg monroe_ionphoton_rtio_core_outputs_gates_record0_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record0_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record0_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record0_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record1_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record1_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record1_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record1_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record2_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record2_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record2_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record2_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record3_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record3_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record3_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record3_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record4_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record4_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record4_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record4_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record5_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record5_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record5_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record5_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record6_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record6_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record6_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record6_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data1 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_gates_record7_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_gates_record7_seqn1 = 12'd0;
wire monroe_ionphoton_rtio_core_outputs_gates_record7_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_gates_record7_nondata_replace_occured;
reg [5:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel1 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address1 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data1 = 32'd0;
wire [60:0] monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp;
reg monroe_ionphoton_rtio_core_outputs_collision = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_collision_channel = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_busy = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_busy_channel = 6'd0;
wire monroe_ionphoton_rtio_core_outputs_record0_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record0_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record0_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record0_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record0_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record0_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record1_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record1_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record1_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record1_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record1_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record1_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record2_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record2_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record2_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record2_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record2_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record2_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record3_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record3_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record3_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record3_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record3_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record3_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record4_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record4_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record4_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record4_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record4_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record4_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record5_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record5_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record5_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record5_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record5_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record5_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record6_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record6_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record6_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record6_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record6_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record6_payload_data2;
wire monroe_ionphoton_rtio_core_outputs_record7_valid0;
wire [11:0] monroe_ionphoton_rtio_core_outputs_record7_seqn2;
wire monroe_ionphoton_rtio_core_outputs_record7_replace_occured;
wire monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured;
wire [5:0] monroe_ionphoton_rtio_core_outputs_record7_payload_channel2;
wire [2:0] monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0;
wire [1:0] monroe_ionphoton_rtio_core_outputs_record7_payload_address2;
wire [31:0] monroe_ionphoton_rtio_core_outputs_record7_payload_data2;
reg monroe_ionphoton_rtio_core_outputs_record0_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record0_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record1_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record1_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record2_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record2_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record3_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record3_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record4_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record4_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record5_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record5_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record6_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record6_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record7_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record7_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference1;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference2;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference3;
reg monroe_ionphoton_rtio_core_outputs_record8_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record8_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record9_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record9_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record10_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record10_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record11_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record11_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record12_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record12_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record13_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record13_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record14_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record14_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record15_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record15_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference4;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference5;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference6;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference7;
reg monroe_ionphoton_rtio_core_outputs_record16_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record16_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record17_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record17_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record18_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record18_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record19_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record19_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record20_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record20_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record21_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record21_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record22_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record22_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record23_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record23_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference8;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference9;
reg monroe_ionphoton_rtio_core_outputs_record24_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record24_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record25_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record25_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record26_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record26_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record27_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record27_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record28_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record28_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record29_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record29_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record30_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record30_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record31_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record31_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference10;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference11;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference12;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference13;
reg monroe_ionphoton_rtio_core_outputs_record32_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record32_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record32_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record32_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record32_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record32_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record32_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record32_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record33_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record33_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record34_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record34_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record35_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record35_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record36_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record36_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record37_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record37_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record38_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record38_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record39_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record39_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record39_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record39_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record39_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record39_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record39_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record39_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference14;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference15;
reg monroe_ionphoton_rtio_core_outputs_record40_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record40_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record40_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record40_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record40_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record40_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record40_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record40_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record41_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record41_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record42_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record42_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record43_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record43_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record44_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record44_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record45_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record45_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record46_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record46_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record47_rec_valid = 1'd0;
reg [11:0] monroe_ionphoton_rtio_core_outputs_record47_rec_seqn = 12'd0;
reg monroe_ionphoton_rtio_core_outputs_record47_rec_replace_occured = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_record47_rec_nondata_replace_occured = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record47_rec_payload_channel = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record47_rec_payload_fine_ts = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record47_rec_payload_address = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record47_rec_payload_data = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference16;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference17;
reg monroe_ionphoton_rtio_core_outputs_nondata_difference18;
reg monroe_ionphoton_rtio_core_outputs_record0_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record0_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record0_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record0_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record1_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record1_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record1_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record1_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record2_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record2_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record2_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record2_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record3_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record3_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record3_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record3_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record4_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record4_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record4_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record4_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record5_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record5_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record5_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record5_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record6_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record6_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record6_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record6_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_record7_valid1 = 1'd0;
wire monroe_ionphoton_rtio_core_outputs_record7_collision;
reg [5:0] monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 = 6'd0;
reg [2:0] monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1 = 3'd0;
reg [1:0] monroe_ionphoton_rtio_core_outputs_record7_payload_address3 = 2'd0;
reg [31:0] monroe_ionphoton_rtio_core_outputs_record7_payload_data3 = 32'd0;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r0 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r0 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory0_adr;
wire monroe_ionphoton_rtio_core_outputs_memory0_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r1 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r1 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory1_adr;
wire monroe_ionphoton_rtio_core_outputs_memory1_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r2 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r2 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory2_adr;
wire monroe_ionphoton_rtio_core_outputs_memory2_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r3 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r3 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory3_adr;
wire monroe_ionphoton_rtio_core_outputs_memory3_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r4 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r4 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory4_adr;
wire monroe_ionphoton_rtio_core_outputs_memory4_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r5 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r5 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory5_adr;
wire monroe_ionphoton_rtio_core_outputs_memory5_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r6 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r6 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory6_adr;
wire monroe_ionphoton_rtio_core_outputs_memory6_dat_r;
reg monroe_ionphoton_rtio_core_outputs_replace_occured_r7 = 1'd0;
reg monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r7 = 1'd0;
wire [5:0] monroe_ionphoton_rtio_core_outputs_memory7_adr;
wire monroe_ionphoton_rtio_core_outputs_memory7_dat_r;
wire monroe_ionphoton_rtio_core_outputs_selected0;
wire monroe_ionphoton_rtio_core_outputs_selected1;
wire monroe_ionphoton_rtio_core_outputs_selected2;
wire monroe_ionphoton_rtio_core_outputs_selected3;
wire monroe_ionphoton_rtio_core_outputs_selected4;
wire monroe_ionphoton_rtio_core_outputs_selected5;
wire monroe_ionphoton_rtio_core_outputs_selected6;
wire monroe_ionphoton_rtio_core_outputs_selected7;
wire monroe_ionphoton_rtio_core_outputs_selected8;
wire monroe_ionphoton_rtio_core_outputs_selected9;
wire monroe_ionphoton_rtio_core_outputs_selected10;
wire monroe_ionphoton_rtio_core_outputs_selected11;
wire monroe_ionphoton_rtio_core_outputs_selected12;
wire monroe_ionphoton_rtio_core_outputs_selected13;
wire monroe_ionphoton_rtio_core_outputs_selected14;
wire monroe_ionphoton_rtio_core_outputs_selected15;
wire monroe_ionphoton_rtio_core_outputs_selected16;
wire monroe_ionphoton_rtio_core_outputs_selected17;
wire monroe_ionphoton_rtio_core_outputs_selected18;
wire monroe_ionphoton_rtio_core_outputs_selected19;
wire monroe_ionphoton_rtio_core_outputs_selected20;
wire monroe_ionphoton_rtio_core_outputs_selected21;
wire monroe_ionphoton_rtio_core_outputs_selected22;
wire monroe_ionphoton_rtio_core_outputs_selected23;
wire monroe_ionphoton_rtio_core_outputs_selected24;
wire monroe_ionphoton_rtio_core_outputs_selected25;
wire monroe_ionphoton_rtio_core_outputs_selected26;
wire monroe_ionphoton_rtio_core_outputs_selected27;
wire monroe_ionphoton_rtio_core_outputs_selected28;
wire monroe_ionphoton_rtio_core_outputs_selected29;
wire monroe_ionphoton_rtio_core_outputs_selected30;
wire monroe_ionphoton_rtio_core_outputs_selected31;
wire monroe_ionphoton_rtio_core_outputs_selected32;
wire monroe_ionphoton_rtio_core_outputs_selected33;
wire monroe_ionphoton_rtio_core_outputs_selected34;
wire monroe_ionphoton_rtio_core_outputs_selected35;
wire monroe_ionphoton_rtio_core_outputs_selected36;
wire monroe_ionphoton_rtio_core_outputs_selected37;
wire monroe_ionphoton_rtio_core_outputs_selected38;
wire monroe_ionphoton_rtio_core_outputs_selected39;
wire monroe_ionphoton_rtio_core_outputs_selected40;
wire monroe_ionphoton_rtio_core_outputs_selected41;
wire monroe_ionphoton_rtio_core_outputs_selected42;
wire monroe_ionphoton_rtio_core_outputs_selected43;
wire monroe_ionphoton_rtio_core_outputs_selected44;
wire monroe_ionphoton_rtio_core_outputs_selected45;
wire monroe_ionphoton_rtio_core_outputs_selected46;
wire monroe_ionphoton_rtio_core_outputs_selected47;
wire monroe_ionphoton_rtio_core_outputs_selected48;
wire monroe_ionphoton_rtio_core_outputs_selected49;
wire monroe_ionphoton_rtio_core_outputs_selected50;
wire monroe_ionphoton_rtio_core_outputs_selected51;
wire monroe_ionphoton_rtio_core_outputs_selected52;
wire monroe_ionphoton_rtio_core_outputs_selected53;
wire monroe_ionphoton_rtio_core_outputs_selected54;
wire monroe_ionphoton_rtio_core_outputs_selected55;
wire monroe_ionphoton_rtio_core_outputs_selected56;
wire monroe_ionphoton_rtio_core_outputs_selected57;
wire monroe_ionphoton_rtio_core_outputs_selected58;
wire monroe_ionphoton_rtio_core_outputs_selected59;
wire monroe_ionphoton_rtio_core_outputs_selected60;
wire monroe_ionphoton_rtio_core_outputs_selected61;
wire monroe_ionphoton_rtio_core_outputs_selected62;
wire monroe_ionphoton_rtio_core_outputs_selected63;
wire monroe_ionphoton_rtio_core_outputs_selected64;
wire monroe_ionphoton_rtio_core_outputs_selected65;
wire monroe_ionphoton_rtio_core_outputs_selected66;
wire monroe_ionphoton_rtio_core_outputs_selected67;
wire monroe_ionphoton_rtio_core_outputs_selected68;
wire monroe_ionphoton_rtio_core_outputs_selected69;
wire monroe_ionphoton_rtio_core_outputs_selected70;
wire monroe_ionphoton_rtio_core_outputs_selected71;
wire monroe_ionphoton_rtio_core_outputs_selected72;
wire monroe_ionphoton_rtio_core_outputs_selected73;
wire monroe_ionphoton_rtio_core_outputs_selected74;
wire monroe_ionphoton_rtio_core_outputs_selected75;
wire monroe_ionphoton_rtio_core_outputs_selected76;
wire monroe_ionphoton_rtio_core_outputs_selected77;
wire monroe_ionphoton_rtio_core_outputs_selected78;
wire monroe_ionphoton_rtio_core_outputs_selected79;
wire monroe_ionphoton_rtio_core_outputs_selected80;
wire monroe_ionphoton_rtio_core_outputs_selected81;
wire monroe_ionphoton_rtio_core_outputs_selected82;
wire monroe_ionphoton_rtio_core_outputs_selected83;
wire monroe_ionphoton_rtio_core_outputs_selected84;
wire monroe_ionphoton_rtio_core_outputs_selected85;
wire monroe_ionphoton_rtio_core_outputs_selected86;
wire monroe_ionphoton_rtio_core_outputs_selected87;
wire monroe_ionphoton_rtio_core_outputs_selected88;
wire monroe_ionphoton_rtio_core_outputs_selected89;
wire monroe_ionphoton_rtio_core_outputs_selected90;
wire monroe_ionphoton_rtio_core_outputs_selected91;
wire monroe_ionphoton_rtio_core_outputs_selected92;
wire monroe_ionphoton_rtio_core_outputs_selected93;
wire monroe_ionphoton_rtio_core_outputs_selected94;
wire monroe_ionphoton_rtio_core_outputs_selected95;
wire monroe_ionphoton_rtio_core_outputs_selected96;
wire monroe_ionphoton_rtio_core_outputs_selected97;
wire monroe_ionphoton_rtio_core_outputs_selected98;
wire monroe_ionphoton_rtio_core_outputs_selected99;
wire monroe_ionphoton_rtio_core_outputs_selected100;
wire monroe_ionphoton_rtio_core_outputs_selected101;
wire monroe_ionphoton_rtio_core_outputs_selected102;
wire monroe_ionphoton_rtio_core_outputs_selected103;
wire monroe_ionphoton_rtio_core_outputs_selected104;
wire monroe_ionphoton_rtio_core_outputs_selected105;
wire monroe_ionphoton_rtio_core_outputs_selected106;
wire monroe_ionphoton_rtio_core_outputs_selected107;
wire monroe_ionphoton_rtio_core_outputs_selected108;
wire monroe_ionphoton_rtio_core_outputs_selected109;
wire monroe_ionphoton_rtio_core_outputs_selected110;
wire monroe_ionphoton_rtio_core_outputs_selected111;
wire monroe_ionphoton_rtio_core_outputs_selected112;
wire monroe_ionphoton_rtio_core_outputs_selected113;
wire monroe_ionphoton_rtio_core_outputs_selected114;
wire monroe_ionphoton_rtio_core_outputs_selected115;
wire monroe_ionphoton_rtio_core_outputs_selected116;
wire monroe_ionphoton_rtio_core_outputs_selected117;
wire monroe_ionphoton_rtio_core_outputs_selected118;
wire monroe_ionphoton_rtio_core_outputs_selected119;
wire monroe_ionphoton_rtio_core_outputs_selected120;
wire monroe_ionphoton_rtio_core_outputs_selected121;
wire monroe_ionphoton_rtio_core_outputs_selected122;
wire monroe_ionphoton_rtio_core_outputs_selected123;
wire monroe_ionphoton_rtio_core_outputs_selected124;
wire monroe_ionphoton_rtio_core_outputs_selected125;
wire monroe_ionphoton_rtio_core_outputs_selected126;
wire monroe_ionphoton_rtio_core_outputs_selected127;
wire monroe_ionphoton_rtio_core_outputs_selected128;
wire monroe_ionphoton_rtio_core_outputs_selected129;
wire monroe_ionphoton_rtio_core_outputs_selected130;
wire monroe_ionphoton_rtio_core_outputs_selected131;
wire monroe_ionphoton_rtio_core_outputs_selected132;
wire monroe_ionphoton_rtio_core_outputs_selected133;
wire monroe_ionphoton_rtio_core_outputs_selected134;
wire monroe_ionphoton_rtio_core_outputs_selected135;
wire monroe_ionphoton_rtio_core_outputs_selected136;
wire monroe_ionphoton_rtio_core_outputs_selected137;
wire monroe_ionphoton_rtio_core_outputs_selected138;
wire monroe_ionphoton_rtio_core_outputs_selected139;
wire monroe_ionphoton_rtio_core_outputs_selected140;
wire monroe_ionphoton_rtio_core_outputs_selected141;
wire monroe_ionphoton_rtio_core_outputs_selected142;
wire monroe_ionphoton_rtio_core_outputs_selected143;
wire monroe_ionphoton_rtio_core_outputs_selected144;
wire monroe_ionphoton_rtio_core_outputs_selected145;
wire monroe_ionphoton_rtio_core_outputs_selected146;
wire monroe_ionphoton_rtio_core_outputs_selected147;
wire monroe_ionphoton_rtio_core_outputs_selected148;
wire monroe_ionphoton_rtio_core_outputs_selected149;
wire monroe_ionphoton_rtio_core_outputs_selected150;
wire monroe_ionphoton_rtio_core_outputs_selected151;
wire monroe_ionphoton_rtio_core_outputs_selected152;
wire monroe_ionphoton_rtio_core_outputs_selected153;
wire monroe_ionphoton_rtio_core_outputs_selected154;
wire monroe_ionphoton_rtio_core_outputs_selected155;
wire monroe_ionphoton_rtio_core_outputs_selected156;
wire monroe_ionphoton_rtio_core_outputs_selected157;
wire monroe_ionphoton_rtio_core_outputs_selected158;
wire monroe_ionphoton_rtio_core_outputs_selected159;
wire monroe_ionphoton_rtio_core_outputs_selected160;
wire monroe_ionphoton_rtio_core_outputs_selected161;
wire monroe_ionphoton_rtio_core_outputs_selected162;
wire monroe_ionphoton_rtio_core_outputs_selected163;
wire monroe_ionphoton_rtio_core_outputs_selected164;
wire monroe_ionphoton_rtio_core_outputs_selected165;
wire monroe_ionphoton_rtio_core_outputs_selected166;
wire monroe_ionphoton_rtio_core_outputs_selected167;
wire monroe_ionphoton_rtio_core_outputs_selected168;
wire monroe_ionphoton_rtio_core_outputs_selected169;
wire monroe_ionphoton_rtio_core_outputs_selected170;
wire monroe_ionphoton_rtio_core_outputs_selected171;
wire monroe_ionphoton_rtio_core_outputs_selected172;
wire monroe_ionphoton_rtio_core_outputs_selected173;
wire monroe_ionphoton_rtio_core_outputs_selected174;
wire monroe_ionphoton_rtio_core_outputs_selected175;
wire monroe_ionphoton_rtio_core_outputs_selected176;
wire monroe_ionphoton_rtio_core_outputs_selected177;
wire monroe_ionphoton_rtio_core_outputs_selected178;
wire monroe_ionphoton_rtio_core_outputs_selected179;
wire monroe_ionphoton_rtio_core_outputs_selected180;
wire monroe_ionphoton_rtio_core_outputs_selected181;
wire monroe_ionphoton_rtio_core_outputs_selected182;
wire monroe_ionphoton_rtio_core_outputs_selected183;
wire monroe_ionphoton_rtio_core_outputs_selected184;
wire monroe_ionphoton_rtio_core_outputs_selected185;
wire monroe_ionphoton_rtio_core_outputs_selected186;
wire monroe_ionphoton_rtio_core_outputs_selected187;
wire monroe_ionphoton_rtio_core_outputs_selected188;
wire monroe_ionphoton_rtio_core_outputs_selected189;
wire monroe_ionphoton_rtio_core_outputs_selected190;
wire monroe_ionphoton_rtio_core_outputs_selected191;
wire monroe_ionphoton_rtio_core_outputs_selected192;
wire monroe_ionphoton_rtio_core_outputs_selected193;
wire monroe_ionphoton_rtio_core_outputs_selected194;
wire monroe_ionphoton_rtio_core_outputs_selected195;
wire monroe_ionphoton_rtio_core_outputs_selected196;
wire monroe_ionphoton_rtio_core_outputs_selected197;
wire monroe_ionphoton_rtio_core_outputs_selected198;
wire monroe_ionphoton_rtio_core_outputs_selected199;
wire monroe_ionphoton_rtio_core_outputs_selected200;
wire monroe_ionphoton_rtio_core_outputs_selected201;
wire monroe_ionphoton_rtio_core_outputs_selected202;
wire monroe_ionphoton_rtio_core_outputs_selected203;
wire monroe_ionphoton_rtio_core_outputs_selected204;
wire monroe_ionphoton_rtio_core_outputs_selected205;
wire monroe_ionphoton_rtio_core_outputs_selected206;
wire monroe_ionphoton_rtio_core_outputs_selected207;
wire monroe_ionphoton_rtio_core_outputs_selected208;
wire monroe_ionphoton_rtio_core_outputs_selected209;
wire monroe_ionphoton_rtio_core_outputs_selected210;
wire monroe_ionphoton_rtio_core_outputs_selected211;
wire monroe_ionphoton_rtio_core_outputs_selected212;
wire monroe_ionphoton_rtio_core_outputs_selected213;
wire monroe_ionphoton_rtio_core_outputs_selected214;
wire monroe_ionphoton_rtio_core_outputs_selected215;
wire monroe_ionphoton_rtio_core_outputs_selected216;
wire monroe_ionphoton_rtio_core_outputs_selected217;
wire monroe_ionphoton_rtio_core_outputs_selected218;
wire monroe_ionphoton_rtio_core_outputs_selected219;
wire monroe_ionphoton_rtio_core_outputs_selected220;
wire monroe_ionphoton_rtio_core_outputs_selected221;
wire monroe_ionphoton_rtio_core_outputs_selected222;
wire monroe_ionphoton_rtio_core_outputs_selected223;
wire monroe_ionphoton_rtio_core_outputs_selected224;
wire monroe_ionphoton_rtio_core_outputs_selected225;
wire monroe_ionphoton_rtio_core_outputs_selected226;
wire monroe_ionphoton_rtio_core_outputs_selected227;
wire monroe_ionphoton_rtio_core_outputs_selected228;
wire monroe_ionphoton_rtio_core_outputs_selected229;
wire monroe_ionphoton_rtio_core_outputs_selected230;
wire monroe_ionphoton_rtio_core_outputs_selected231;
wire monroe_ionphoton_rtio_core_outputs_selected232;
wire monroe_ionphoton_rtio_core_outputs_selected233;
wire monroe_ionphoton_rtio_core_outputs_selected234;
wire monroe_ionphoton_rtio_core_outputs_selected235;
wire monroe_ionphoton_rtio_core_outputs_selected236;
wire monroe_ionphoton_rtio_core_outputs_selected237;
wire monroe_ionphoton_rtio_core_outputs_selected238;
wire monroe_ionphoton_rtio_core_outputs_selected239;
wire monroe_ionphoton_rtio_core_outputs_selected240;
wire monroe_ionphoton_rtio_core_outputs_selected241;
wire monroe_ionphoton_rtio_core_outputs_selected242;
wire monroe_ionphoton_rtio_core_outputs_selected243;
wire monroe_ionphoton_rtio_core_outputs_selected244;
wire monroe_ionphoton_rtio_core_outputs_selected245;
wire monroe_ionphoton_rtio_core_outputs_selected246;
wire monroe_ionphoton_rtio_core_outputs_selected247;
wire monroe_ionphoton_rtio_core_outputs_selected248;
wire monroe_ionphoton_rtio_core_outputs_selected249;
wire monroe_ionphoton_rtio_core_outputs_selected250;
wire monroe_ionphoton_rtio_core_outputs_selected251;
wire monroe_ionphoton_rtio_core_outputs_selected252;
wire monroe_ionphoton_rtio_core_outputs_selected253;
wire monroe_ionphoton_rtio_core_outputs_selected254;
wire monroe_ionphoton_rtio_core_outputs_selected255;
wire monroe_ionphoton_rtio_core_outputs_selected256;
wire monroe_ionphoton_rtio_core_outputs_selected257;
wire monroe_ionphoton_rtio_core_outputs_selected258;
wire monroe_ionphoton_rtio_core_outputs_selected259;
wire monroe_ionphoton_rtio_core_outputs_selected260;
wire monroe_ionphoton_rtio_core_outputs_selected261;
wire monroe_ionphoton_rtio_core_outputs_selected262;
wire monroe_ionphoton_rtio_core_outputs_selected263;
wire monroe_ionphoton_rtio_core_outputs_selected264;
wire monroe_ionphoton_rtio_core_outputs_selected265;
wire monroe_ionphoton_rtio_core_outputs_selected266;
wire monroe_ionphoton_rtio_core_outputs_selected267;
wire monroe_ionphoton_rtio_core_outputs_selected268;
wire monroe_ionphoton_rtio_core_outputs_selected269;
wire monroe_ionphoton_rtio_core_outputs_selected270;
wire monroe_ionphoton_rtio_core_outputs_selected271;
wire monroe_ionphoton_rtio_core_outputs_selected272;
wire monroe_ionphoton_rtio_core_outputs_selected273;
wire monroe_ionphoton_rtio_core_outputs_selected274;
wire monroe_ionphoton_rtio_core_outputs_selected275;
wire monroe_ionphoton_rtio_core_outputs_selected276;
wire monroe_ionphoton_rtio_core_outputs_selected277;
wire monroe_ionphoton_rtio_core_outputs_selected278;
wire monroe_ionphoton_rtio_core_outputs_selected279;
wire monroe_ionphoton_rtio_core_outputs_selected280;
wire monroe_ionphoton_rtio_core_outputs_selected281;
wire monroe_ionphoton_rtio_core_outputs_selected282;
wire monroe_ionphoton_rtio_core_outputs_selected283;
wire monroe_ionphoton_rtio_core_outputs_selected284;
wire monroe_ionphoton_rtio_core_outputs_selected285;
wire monroe_ionphoton_rtio_core_outputs_selected286;
wire monroe_ionphoton_rtio_core_outputs_selected287;
wire monroe_ionphoton_rtio_core_outputs_selected288;
wire monroe_ionphoton_rtio_core_outputs_selected289;
wire monroe_ionphoton_rtio_core_outputs_selected290;
wire monroe_ionphoton_rtio_core_outputs_selected291;
wire monroe_ionphoton_rtio_core_outputs_selected292;
wire monroe_ionphoton_rtio_core_outputs_selected293;
wire monroe_ionphoton_rtio_core_outputs_selected294;
wire monroe_ionphoton_rtio_core_outputs_selected295;
reg monroe_ionphoton_rtio_core_outputs_stb_r0 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r0 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r1 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r1 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r2 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r2 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r3 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r3 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r4 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r4 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r5 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r5 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r6 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r6 = 6'd0;
reg monroe_ionphoton_rtio_core_outputs_stb_r7 = 1'd0;
reg [5:0] monroe_ionphoton_rtio_core_outputs_channel_r7 = 6'd0;
reg monroe_ionphoton_rtio_core_inputs_i_ack = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_readable;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_produce_rdomain;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_consume_wdomain;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_we;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_dat_w;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_record0_fifo_in_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record0_fifo_in_timestamp;
wire monroe_ionphoton_rtio_core_inputs_record0_fifo_out_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record0_fifo_out_timestamp;
wire monroe_ionphoton_rtio_core_inputs_overflow_io0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer0_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected0;
reg monroe_ionphoton_rtio_core_inputs_overflow0 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_readable;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_produce_rdomain;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_consume_wdomain;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_we;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_dat_w;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_record1_fifo_in_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record1_fifo_in_timestamp;
wire monroe_ionphoton_rtio_core_inputs_record1_fifo_out_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record1_fifo_out_timestamp;
wire monroe_ionphoton_rtio_core_inputs_overflow_io1;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer1_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected1;
reg monroe_ionphoton_rtio_core_inputs_overflow1 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_readable;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_produce_rdomain;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_consume_wdomain;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_we;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_dat_w;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_record2_fifo_in_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record2_fifo_in_timestamp;
wire monroe_ionphoton_rtio_core_inputs_record2_fifo_out_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record2_fifo_out_timestamp;
wire monroe_ionphoton_rtio_core_inputs_overflow_io2;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer2_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected2;
reg monroe_ionphoton_rtio_core_inputs_overflow2 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_readable;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_ce;
(* dont_touch = "true" *) reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q = 7'd0;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_binary = 7'd0;
reg [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_produce_rdomain;
wire [6:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_consume_wdomain;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_we;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_dat_w;
wire [5:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_adr;
wire [64:0] monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_record3_fifo_in_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record3_fifo_in_timestamp;
wire monroe_ionphoton_rtio_core_inputs_record3_fifo_out_data;
wire [63:0] monroe_ionphoton_rtio_core_inputs_record3_fifo_out_timestamp;
wire monroe_ionphoton_rtio_core_inputs_overflow_io3;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer3_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected3;
reg monroe_ionphoton_rtio_core_inputs_overflow3 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_readable;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_produce_rdomain;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_consume_wdomain;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_we;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_dat_w;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_dat_r;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record4_fifo_in_data;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record4_fifo_out_data;
wire monroe_ionphoton_rtio_core_inputs_overflow_io4;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer4_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected4;
reg monroe_ionphoton_rtio_core_inputs_overflow4 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_readable;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_produce_rdomain;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_consume_wdomain;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_we;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_dat_w;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_dat_r;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record5_fifo_in_data;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record5_fifo_out_data;
wire monroe_ionphoton_rtio_core_inputs_overflow_io5;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer5_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected5;
reg monroe_ionphoton_rtio_core_inputs_overflow5 = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_we;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_writable;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_re;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_readable;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_ce;
(* dont_touch = "true" *) reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q = 3'd0;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_binary = 3'd0;
reg [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_produce_rdomain;
wire [2:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_consume_wdomain;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_dat_r;
wire monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_we;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_dat_w;
wire [1:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_adr;
wire [31:0] monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_dat_r;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record6_fifo_in_data;
wire [31:0] monroe_ionphoton_rtio_core_inputs_record6_fifo_out_data;
wire monroe_ionphoton_rtio_core_inputs_overflow_io6;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_o;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_i;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_inputs_blindtransfer6_blind = 1'd0;
wire monroe_ionphoton_rtio_core_inputs_selected6;
reg monroe_ionphoton_rtio_core_inputs_overflow6 = 1'd0;
wire [1:0] monroe_ionphoton_rtio_core_inputs_i_status_raw;
reg [63:0] monroe_ionphoton_rtio_core_inputs_input_timeout = 64'd0;
reg monroe_ionphoton_rtio_core_inputs_input_pending = 1'd0;
wire monroe_ionphoton_rtio_core_o_collision_sync_i;
wire monroe_ionphoton_rtio_core_o_collision_sync_o;
wire [15:0] monroe_ionphoton_rtio_core_o_collision_sync_data_i;
wire [15:0] monroe_ionphoton_rtio_core_o_collision_sync_data_o;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_i;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_o;
reg monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o;
reg monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_i;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_o;
reg monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_o_collision_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] monroe_ionphoton_rtio_core_o_collision_sync_bxfer_data = 16'd0;
wire monroe_ionphoton_rtio_core_o_busy_sync_i;
wire monroe_ionphoton_rtio_core_o_busy_sync_o;
wire [15:0] monroe_ionphoton_rtio_core_o_busy_sync_data_i;
wire [15:0] monroe_ionphoton_rtio_core_o_busy_sync_data_o;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_i;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_o;
reg monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o;
reg monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o_r = 1'd0;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_i;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_o;
reg monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_i = 1'd0;
wire monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o;
reg monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o_r = 1'd0;
reg monroe_ionphoton_rtio_core_o_busy_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] monroe_ionphoton_rtio_core_o_busy_sync_bxfer_data = 16'd0;
reg monroe_ionphoton_rtio_core_o_collision = 1'd0;
reg monroe_ionphoton_rtio_core_o_busy = 1'd0;
reg monroe_ionphoton_rtio_core_o_sequence_error = 1'd0;
reg [31:0] monroe_ionphoton_rtio_target_storage_full = 32'd0;
wire [31:0] monroe_ionphoton_rtio_target_storage;
reg monroe_ionphoton_rtio_target_re = 1'd0;
wire monroe_ionphoton_rtio_now_hi_re;
wire [31:0] monroe_ionphoton_rtio_now_hi_r;
wire [31:0] monroe_ionphoton_rtio_now_hi_w;
wire monroe_ionphoton_rtio_now_lo_re;
wire [31:0] monroe_ionphoton_rtio_now_lo_r;
wire [31:0] monroe_ionphoton_rtio_now_lo_w;
reg [511:0] monroe_ionphoton_rtio_o_data_storage_full = 512'd0;
wire [511:0] monroe_ionphoton_rtio_o_data_storage;
reg monroe_ionphoton_rtio_o_data_re = 1'd0;
wire monroe_ionphoton_rtio_o_data_we;
wire [511:0] monroe_ionphoton_rtio_o_data_dat_w;
wire [2:0] monroe_ionphoton_rtio_o_status_status;
reg [63:0] monroe_ionphoton_rtio_i_timeout_storage_full = 64'd0;
wire [63:0] monroe_ionphoton_rtio_i_timeout_storage;
reg monroe_ionphoton_rtio_i_timeout_re = 1'd0;
wire [31:0] monroe_ionphoton_rtio_i_data_status;
wire [63:0] monroe_ionphoton_rtio_i_timestamp_status;
wire [3:0] monroe_ionphoton_rtio_i_status_status;
wire monroe_ionphoton_rtio_i_overflow_reset_re;
wire monroe_ionphoton_rtio_i_overflow_reset_r;
reg monroe_ionphoton_rtio_i_overflow_reset_w = 1'd0;
reg [63:0] monroe_ionphoton_rtio_counter_status = 64'd0;
wire monroe_ionphoton_rtio_counter_update_re;
wire monroe_ionphoton_rtio_counter_update_r;
reg monroe_ionphoton_rtio_counter_update_w = 1'd0;
reg [1:0] monroe_ionphoton_rtio_cri_cmd;
wire [23:0] monroe_ionphoton_rtio_cri_chan_sel;
wire [63:0] monroe_ionphoton_rtio_cri_o_timestamp;
wire [511:0] monroe_ionphoton_rtio_cri_o_data;
wire [7:0] monroe_ionphoton_rtio_cri_o_address;
wire [2:0] monroe_ionphoton_rtio_cri_o_status;
wire monroe_ionphoton_rtio_cri_o_buffer_space_valid;
wire [15:0] monroe_ionphoton_rtio_cri_o_buffer_space;
wire [63:0] monroe_ionphoton_rtio_cri_i_timeout;
wire [31:0] monroe_ionphoton_rtio_cri_i_data;
wire [63:0] monroe_ionphoton_rtio_cri_i_timestamp;
wire [3:0] monroe_ionphoton_rtio_cri_i_status;
reg [31:0] monroe_ionphoton_rtio_now_hi_backing = 32'd0;
reg [63:0] monroe_ionphoton_rtio_now = 64'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_adr;
reg [127:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_dat_w = 128'd0;
wire [127:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_dat_r;
reg [15:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_sel = 16'd0;
wire monroe_ionphoton_monroe_ionphoton_interface0_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_interface0_bus_stb;
wire monroe_ionphoton_monroe_ionphoton_interface0_bus_ack;
reg monroe_ionphoton_monroe_ionphoton_interface0_bus_we = 1'd0;
reg [2:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_cti = 3'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_interface0_bus_bte = 2'd0;
wire monroe_ionphoton_monroe_ionphoton_interface0_bus_err;
wire monroe_ionphoton_dma_enable_enable_re;
wire monroe_ionphoton_dma_enable_enable_r;
reg monroe_ionphoton_dma_enable_enable_w;
reg monroe_ionphoton_dma_flow_enable;
reg monroe_ionphoton_dma_dma_sink_stb = 1'd0;
wire monroe_ionphoton_dma_dma_sink_ack;
reg monroe_ionphoton_dma_dma_sink_eop = 1'd0;
reg [29:0] monroe_ionphoton_dma_dma_sink_payload_address = 30'd0;
wire monroe_ionphoton_dma_dma_source_stb;
wire monroe_ionphoton_dma_dma_source_ack;
reg monroe_ionphoton_dma_dma_source_eop = 1'd0;
reg [127:0] monroe_ionphoton_dma_dma_source_payload_data = 128'd0;
wire monroe_ionphoton_dma_dma_bus_stb;
reg monroe_ionphoton_dma_dma_data_reg_loaded = 1'd0;
reg [33:0] monroe_ionphoton_dma_dma_storage_full = 34'd0;
wire [29:0] monroe_ionphoton_dma_dma_storage;
reg monroe_ionphoton_dma_dma_re = 1'd0;
reg monroe_ionphoton_dma_dma_enable_r = 1'd0;
wire monroe_ionphoton_dma_rawslicer_sink_stb;
reg monroe_ionphoton_dma_rawslicer_sink_ack;
wire monroe_ionphoton_dma_rawslicer_sink_eop;
wire [127:0] monroe_ionphoton_dma_rawslicer_sink_payload_data;
wire [615:0] monroe_ionphoton_dma_rawslicer_source;
reg monroe_ionphoton_dma_rawslicer_source_stb;
reg [6:0] monroe_ionphoton_dma_rawslicer_source_consume;
reg monroe_ionphoton_dma_rawslicer_flush;
reg monroe_ionphoton_dma_rawslicer_flush_done;
reg [735:0] monroe_ionphoton_dma_rawslicer_buf = 736'd0;
reg [6:0] monroe_ionphoton_dma_rawslicer_level = 7'd0;
reg [6:0] monroe_ionphoton_dma_rawslicer_next_level;
reg monroe_ionphoton_dma_rawslicer_load_buf;
reg monroe_ionphoton_dma_rawslicer_shift_buf;
reg monroe_ionphoton_dma_reset = 1'd0;
reg monroe_ionphoton_dma_record_converter_source_stb;
wire monroe_ionphoton_dma_record_converter_source_ack;
reg monroe_ionphoton_dma_record_converter_source_eop;
reg [7:0] monroe_ionphoton_dma_record_converter_source_payload_length = 8'd0;
wire [23:0] monroe_ionphoton_dma_record_converter_source_payload_channel;
wire [63:0] monroe_ionphoton_dma_record_converter_source_payload_timestamp;
wire [7:0] monroe_ionphoton_dma_record_converter_source_payload_address;
reg [511:0] monroe_ionphoton_dma_record_converter_source_payload_data;
reg monroe_ionphoton_dma_record_converter_end_marker_found;
reg monroe_ionphoton_dma_record_converter_flush;
wire [7:0] monroe_ionphoton_dma_record_converter_record_raw_length;
wire [23:0] monroe_ionphoton_dma_record_converter_record_raw_channel;
wire [63:0] monroe_ionphoton_dma_record_converter_record_raw_timestamp;
wire [7:0] monroe_ionphoton_dma_record_converter_record_raw_address;
wire [511:0] monroe_ionphoton_dma_record_converter_record_raw_data;
reg [63:0] monroe_ionphoton_dma_time_offset_storage_full = 64'd0;
wire [63:0] monroe_ionphoton_dma_time_offset_storage;
reg monroe_ionphoton_dma_time_offset_re = 1'd0;
reg monroe_ionphoton_dma_time_offset_source_stb = 1'd0;
wire monroe_ionphoton_dma_time_offset_source_ack;
reg monroe_ionphoton_dma_time_offset_source_eop = 1'd0;
reg [7:0] monroe_ionphoton_dma_time_offset_source_payload_length = 8'd0;
reg [23:0] monroe_ionphoton_dma_time_offset_source_payload_channel = 24'd0;
reg [63:0] monroe_ionphoton_dma_time_offset_source_payload_timestamp = 64'd0;
reg [7:0] monroe_ionphoton_dma_time_offset_source_payload_address = 8'd0;
reg [511:0] monroe_ionphoton_dma_time_offset_source_payload_data = 512'd0;
wire monroe_ionphoton_dma_time_offset_sink_stb;
wire monroe_ionphoton_dma_time_offset_sink_ack;
wire monroe_ionphoton_dma_time_offset_sink_eop;
wire [7:0] monroe_ionphoton_dma_time_offset_sink_payload_length;
wire [23:0] monroe_ionphoton_dma_time_offset_sink_payload_channel;
wire [63:0] monroe_ionphoton_dma_time_offset_sink_payload_timestamp;
wire [7:0] monroe_ionphoton_dma_time_offset_sink_payload_address;
wire [511:0] monroe_ionphoton_dma_time_offset_sink_payload_data;
wire monroe_ionphoton_dma_cri_master_error_re;
wire [1:0] monroe_ionphoton_dma_cri_master_error_r;
reg [1:0] monroe_ionphoton_dma_cri_master_error_w = 2'd0;
reg [23:0] monroe_ionphoton_dma_cri_master_error_channel_status = 24'd0;
reg [63:0] monroe_ionphoton_dma_cri_master_error_timestamp_status = 64'd0;
reg [15:0] monroe_ionphoton_dma_cri_master_error_address_status = 16'd0;
wire monroe_ionphoton_dma_cri_master_sink_stb;
reg monroe_ionphoton_dma_cri_master_sink_ack;
wire monroe_ionphoton_dma_cri_master_sink_eop;
wire [7:0] monroe_ionphoton_dma_cri_master_sink_payload_length;
wire [23:0] monroe_ionphoton_dma_cri_master_sink_payload_channel;
wire [63:0] monroe_ionphoton_dma_cri_master_sink_payload_timestamp;
wire [7:0] monroe_ionphoton_dma_cri_master_sink_payload_address;
wire [511:0] monroe_ionphoton_dma_cri_master_sink_payload_data;
reg [1:0] monroe_ionphoton_dma_cri_master_cri_cmd;
wire [23:0] monroe_ionphoton_dma_cri_master_cri_chan_sel;
wire [63:0] monroe_ionphoton_dma_cri_master_cri_o_timestamp;
wire [511:0] monroe_ionphoton_dma_cri_master_cri_o_data;
wire [7:0] monroe_ionphoton_dma_cri_master_cri_o_address;
wire [2:0] monroe_ionphoton_dma_cri_master_cri_o_status;
wire monroe_ionphoton_dma_cri_master_cri_o_buffer_space_valid;
wire [15:0] monroe_ionphoton_dma_cri_master_cri_o_buffer_space;
reg [63:0] monroe_ionphoton_dma_cri_master_cri_i_timeout = 64'd0;
wire [31:0] monroe_ionphoton_dma_cri_master_cri_i_data;
wire [63:0] monroe_ionphoton_dma_cri_master_cri_i_timestamp;
wire [3:0] monroe_ionphoton_dma_cri_master_cri_i_status;
reg monroe_ionphoton_dma_cri_master_busy;
reg monroe_ionphoton_dma_cri_master_underflow_trigger;
reg monroe_ionphoton_dma_cri_master_link_error_trigger;
wire [29:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank0_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_csrbank0_bus_err = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_target0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_target0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_target0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_re;
wire [2:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_r;
wire [2:0] monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_re;
wire [3:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_r;
wire [3:0] monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_w;
wire [29:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank1_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_csrbank1_bus_err = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_re;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_r;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_re;
wire [23:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_r;
wire [23:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_re;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_r;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_w;
wire monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_re;
wire [15:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_r;
wire [15:0] monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_w;
wire [1:0] monroe_ionphoton_cri_con_shared_cmd;
wire [23:0] monroe_ionphoton_cri_con_shared_chan_sel;
wire [63:0] monroe_ionphoton_cri_con_shared_o_timestamp;
wire [511:0] monroe_ionphoton_cri_con_shared_o_data;
wire [7:0] monroe_ionphoton_cri_con_shared_o_address;
reg [2:0] monroe_ionphoton_cri_con_shared_o_status;
reg monroe_ionphoton_cri_con_shared_o_buffer_space_valid;
reg [15:0] monroe_ionphoton_cri_con_shared_o_buffer_space;
wire [63:0] monroe_ionphoton_cri_con_shared_i_timeout;
reg [31:0] monroe_ionphoton_cri_con_shared_i_data;
reg [63:0] monroe_ionphoton_cri_con_shared_i_timestamp;
reg [3:0] monroe_ionphoton_cri_con_shared_i_status;
reg [1:0] monroe_ionphoton_cri_con_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_cri_con_storage;
reg monroe_ionphoton_cri_con_re = 1'd0;
reg monroe_ionphoton_cri_con_selected = 1'd0;
wire [29:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_adr;
wire [31:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_w;
reg [31:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_r = 32'd0;
wire [3:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_csrbank2_bus_stb;
reg monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank2_bus_we;
wire [2:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cti;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank2_bus_bte;
reg monroe_ionphoton_monroe_ionphoton_csrbank2_bus_err = 1'd0;
wire monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_re;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_r;
wire [1:0] monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_w;
reg [5:0] monroe_ionphoton_mon_chan_sel_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_mon_chan_sel_storage;
reg monroe_ionphoton_mon_chan_sel_re = 1'd0;
reg monroe_ionphoton_mon_probe_sel_storage_full = 1'd0;
wire monroe_ionphoton_mon_probe_sel_storage;
reg monroe_ionphoton_mon_probe_sel_re = 1'd0;
wire monroe_ionphoton_mon_value_update_re;
wire monroe_ionphoton_mon_value_update_r;
reg monroe_ionphoton_mon_value_update_w = 1'd0;
reg monroe_ionphoton_mon_status = 1'd0;
wire monroe_ionphoton_mon_bussynchronizer0_i;
wire monroe_ionphoton_mon_bussynchronizer0_o;
wire monroe_ionphoton_mon_bussynchronizer1_i;
wire monroe_ionphoton_mon_bussynchronizer1_o;
wire monroe_ionphoton_mon_bussynchronizer2_i;
wire monroe_ionphoton_mon_bussynchronizer2_o;
wire monroe_ionphoton_mon_bussynchronizer3_i;
wire monroe_ionphoton_mon_bussynchronizer3_o;
wire monroe_ionphoton_mon_bussynchronizer4_i;
wire monroe_ionphoton_mon_bussynchronizer4_o;
wire monroe_ionphoton_mon_bussynchronizer5_i;
wire monroe_ionphoton_mon_bussynchronizer5_o;
wire monroe_ionphoton_mon_bussynchronizer6_i;
wire monroe_ionphoton_mon_bussynchronizer6_o;
wire monroe_ionphoton_mon_bussynchronizer7_i;
wire monroe_ionphoton_mon_bussynchronizer7_o;
wire monroe_ionphoton_mon_bussynchronizer8_i;
wire monroe_ionphoton_mon_bussynchronizer8_o;
wire monroe_ionphoton_mon_bussynchronizer9_i;
wire monroe_ionphoton_mon_bussynchronizer9_o;
wire monroe_ionphoton_mon_bussynchronizer10_i;
wire monroe_ionphoton_mon_bussynchronizer10_o;
wire monroe_ionphoton_mon_bussynchronizer11_i;
wire monroe_ionphoton_mon_bussynchronizer11_o;
wire monroe_ionphoton_mon_bussynchronizer12_i;
wire monroe_ionphoton_mon_bussynchronizer12_o;
wire monroe_ionphoton_mon_bussynchronizer13_i;
wire monroe_ionphoton_mon_bussynchronizer13_o;
wire monroe_ionphoton_mon_bussynchronizer14_i;
wire monroe_ionphoton_mon_bussynchronizer14_o;
wire monroe_ionphoton_mon_bussynchronizer15_i;
wire monroe_ionphoton_mon_bussynchronizer15_o;
wire monroe_ionphoton_mon_bussynchronizer16_i;
wire monroe_ionphoton_mon_bussynchronizer16_o;
wire monroe_ionphoton_mon_bussynchronizer17_i;
wire monroe_ionphoton_mon_bussynchronizer17_o;
wire monroe_ionphoton_mon_bussynchronizer18_i;
wire monroe_ionphoton_mon_bussynchronizer18_o;
wire monroe_ionphoton_mon_bussynchronizer19_i;
wire monroe_ionphoton_mon_bussynchronizer19_o;
wire monroe_ionphoton_mon_bussynchronizer20_i;
wire monroe_ionphoton_mon_bussynchronizer20_o;
wire monroe_ionphoton_mon_bussynchronizer21_i;
wire monroe_ionphoton_mon_bussynchronizer21_o;
wire monroe_ionphoton_mon_bussynchronizer22_i;
wire monroe_ionphoton_mon_bussynchronizer22_o;
wire monroe_ionphoton_mon_bussynchronizer23_i;
wire monroe_ionphoton_mon_bussynchronizer23_o;
wire monroe_ionphoton_mon_bussynchronizer24_i;
wire monroe_ionphoton_mon_bussynchronizer24_o;
wire monroe_ionphoton_mon_bussynchronizer25_i;
wire monroe_ionphoton_mon_bussynchronizer25_o;
wire monroe_ionphoton_mon_bussynchronizer26_i;
wire monroe_ionphoton_mon_bussynchronizer26_o;
wire monroe_ionphoton_mon_bussynchronizer27_i;
wire monroe_ionphoton_mon_bussynchronizer27_o;
wire monroe_ionphoton_mon_bussynchronizer28_i;
wire monroe_ionphoton_mon_bussynchronizer28_o;
wire monroe_ionphoton_mon_bussynchronizer29_i;
wire monroe_ionphoton_mon_bussynchronizer29_o;
wire monroe_ionphoton_mon_bussynchronizer30_i;
wire monroe_ionphoton_mon_bussynchronizer30_o;
wire monroe_ionphoton_mon_bussynchronizer31_i;
wire monroe_ionphoton_mon_bussynchronizer31_o;
wire monroe_ionphoton_mon_bussynchronizer32_i;
wire monroe_ionphoton_mon_bussynchronizer32_o;
wire monroe_ionphoton_mon_bussynchronizer33_i;
wire monroe_ionphoton_mon_bussynchronizer33_o;
wire monroe_ionphoton_mon_bussynchronizer34_i;
wire monroe_ionphoton_mon_bussynchronizer34_o;
wire monroe_ionphoton_mon_bussynchronizer35_i;
wire monroe_ionphoton_mon_bussynchronizer35_o;
wire monroe_ionphoton_mon_bussynchronizer36_i;
wire monroe_ionphoton_mon_bussynchronizer36_o;
reg [5:0] monroe_ionphoton_inj_chan_sel_storage_full = 6'd0;
wire [5:0] monroe_ionphoton_inj_chan_sel_storage;
reg monroe_ionphoton_inj_chan_sel_re = 1'd0;
reg [1:0] monroe_ionphoton_inj_override_sel_storage_full = 2'd0;
wire [1:0] monroe_ionphoton_inj_override_sel_storage;
reg monroe_ionphoton_inj_override_sel_re = 1'd0;
wire monroe_ionphoton_inj_value_re;
wire monroe_ionphoton_inj_value_r;
wire monroe_ionphoton_inj_value_w;
reg monroe_ionphoton_inj_o_sys0 = 1'd0;
reg monroe_ionphoton_inj_o_sys1 = 1'd0;
reg monroe_ionphoton_inj_o_sys2 = 1'd0;
reg monroe_ionphoton_inj_o_sys3 = 1'd0;
reg monroe_ionphoton_inj_o_sys4 = 1'd0;
reg monroe_ionphoton_inj_o_sys5 = 1'd0;
reg monroe_ionphoton_inj_o_sys6 = 1'd0;
reg monroe_ionphoton_inj_o_sys7 = 1'd0;
reg monroe_ionphoton_inj_o_sys8 = 1'd0;
reg monroe_ionphoton_inj_o_sys9 = 1'd0;
reg monroe_ionphoton_inj_o_sys10 = 1'd0;
reg monroe_ionphoton_inj_o_sys11 = 1'd0;
reg monroe_ionphoton_inj_o_sys12 = 1'd0;
reg monroe_ionphoton_inj_o_sys13 = 1'd0;
reg monroe_ionphoton_inj_o_sys14 = 1'd0;
reg monroe_ionphoton_inj_o_sys15 = 1'd0;
reg monroe_ionphoton_inj_o_sys16 = 1'd0;
reg monroe_ionphoton_inj_o_sys17 = 1'd0;
reg monroe_ionphoton_inj_o_sys18 = 1'd0;
reg monroe_ionphoton_inj_o_sys19 = 1'd0;
reg monroe_ionphoton_inj_o_sys20 = 1'd0;
reg monroe_ionphoton_inj_o_sys21 = 1'd0;
reg monroe_ionphoton_inj_o_sys22 = 1'd0;
reg monroe_ionphoton_inj_o_sys23 = 1'd0;
reg monroe_ionphoton_inj_o_sys24 = 1'd0;
reg monroe_ionphoton_inj_o_sys25 = 1'd0;
reg monroe_ionphoton_inj_o_sys26 = 1'd0;
reg monroe_ionphoton_inj_o_sys27 = 1'd0;
reg monroe_ionphoton_inj_o_sys28 = 1'd0;
reg monroe_ionphoton_inj_o_sys29 = 1'd0;
reg monroe_ionphoton_inj_o_sys30 = 1'd0;
reg monroe_ionphoton_inj_o_sys31 = 1'd0;
reg monroe_ionphoton_inj_o_sys32 = 1'd0;
reg monroe_ionphoton_inj_o_sys33 = 1'd0;
reg monroe_ionphoton_inj_o_sys34 = 1'd0;
reg monroe_ionphoton_inj_o_sys35 = 1'd0;
reg monroe_ionphoton_inj_o_sys36 = 1'd0;
reg monroe_ionphoton_inj_o_sys37 = 1'd0;
reg monroe_ionphoton_inj_o_sys38 = 1'd0;
reg monroe_ionphoton_inj_o_sys39 = 1'd0;
reg monroe_ionphoton_inj_o_sys40 = 1'd0;
reg monroe_ionphoton_inj_o_sys41 = 1'd0;
reg monroe_ionphoton_inj_o_sys42 = 1'd0;
reg monroe_ionphoton_inj_o_sys43 = 1'd0;
reg monroe_ionphoton_inj_o_sys44 = 1'd0;
reg monroe_ionphoton_inj_o_sys45 = 1'd0;
reg monroe_ionphoton_inj_o_sys46 = 1'd0;
reg monroe_ionphoton_inj_o_sys47 = 1'd0;
reg monroe_ionphoton_inj_o_sys48 = 1'd0;
reg monroe_ionphoton_inj_o_sys49 = 1'd0;
reg monroe_ionphoton_inj_o_sys50 = 1'd0;
reg monroe_ionphoton_inj_o_sys51 = 1'd0;
reg monroe_ionphoton_inj_o_sys52 = 1'd0;
reg monroe_ionphoton_inj_o_sys53 = 1'd0;
reg monroe_ionphoton_inj_o_sys54 = 1'd0;
reg monroe_ionphoton_inj_o_sys55 = 1'd0;
reg monroe_ionphoton_inj_o_sys56 = 1'd0;
reg monroe_ionphoton_inj_o_sys57 = 1'd0;
reg monroe_ionphoton_inj_o_sys58 = 1'd0;
reg monroe_ionphoton_inj_o_sys59 = 1'd0;
reg monroe_ionphoton_inj_o_sys60 = 1'd0;
reg monroe_ionphoton_inj_o_sys61 = 1'd0;
reg monroe_ionphoton_inj_o_sys62 = 1'd0;
reg monroe_ionphoton_inj_o_sys63 = 1'd0;
reg monroe_ionphoton_inj_o_sys64 = 1'd0;
reg monroe_ionphoton_inj_o_sys65 = 1'd0;
reg monroe_ionphoton_inj_o_sys66 = 1'd0;
reg monroe_ionphoton_inj_o_sys67 = 1'd0;
reg monroe_ionphoton_inj_o_sys68 = 1'd0;
reg monroe_ionphoton_inj_o_sys69 = 1'd0;
reg [29:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_adr = 30'd0;
wire [127:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_dat_w;
wire [127:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_dat_r;
wire [15:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_sel;
wire monroe_ionphoton_monroe_ionphoton_interface1_bus_cyc;
wire monroe_ionphoton_monroe_ionphoton_interface1_bus_stb;
wire monroe_ionphoton_monroe_ionphoton_interface1_bus_ack;
wire monroe_ionphoton_monroe_ionphoton_interface1_bus_we;
reg [2:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_cti = 3'd0;
reg [1:0] monroe_ionphoton_monroe_ionphoton_interface1_bus_bte = 2'd0;
wire monroe_ionphoton_monroe_ionphoton_interface1_bus_err;
reg monroe_ionphoton_rtio_analyzer_enable_storage_full = 1'd0;
wire monroe_ionphoton_rtio_analyzer_enable_storage;
reg monroe_ionphoton_rtio_analyzer_enable_re = 1'd0;
reg monroe_ionphoton_rtio_analyzer_busy_status = 1'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_source_stb = 1'd0;
wire monroe_ionphoton_rtio_analyzer_message_encoder_source_ack;
reg monroe_ionphoton_rtio_analyzer_message_encoder_source_eop = 1'd0;
reg [255:0] monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data = 256'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_status = 1'd0;
wire monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_re;
wire monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_r;
reg monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_w = 1'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_read_wait_event_r = 1'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_read_done;
reg monroe_ionphoton_rtio_analyzer_message_encoder_read_overflow;
wire monroe_ionphoton_rtio_analyzer_message_encoder_input_output_stb;
reg [1:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_message_type;
wire [29:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_channel;
reg [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_timestamp;
wire [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_rtio_counter;
wire [31:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_address_padding;
reg [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_input_output_data;
reg monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb;
wire [1:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_message_type;
wire [29:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_channel;
reg [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_padding0 = 64'd0;
wire [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_rtio_counter;
reg [7:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_exception_type;
reg [87:0] monroe_ionphoton_rtio_analyzer_message_encoder_exception_padding1 = 88'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_just_written = 1'd0;
wire [1:0] monroe_ionphoton_rtio_analyzer_message_encoder_stopped_message_type;
reg [93:0] monroe_ionphoton_rtio_analyzer_message_encoder_stopped_padding0 = 94'd0;
wire [63:0] monroe_ionphoton_rtio_analyzer_message_encoder_stopped_rtio_counter;
reg [95:0] monroe_ionphoton_rtio_analyzer_message_encoder_stopped_padding1 = 96'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_enable_r = 1'd0;
reg monroe_ionphoton_rtio_analyzer_message_encoder_stopping = 1'd0;
wire monroe_ionphoton_rtio_analyzer_fifo_sink_stb;
wire monroe_ionphoton_rtio_analyzer_fifo_sink_ack;
wire monroe_ionphoton_rtio_analyzer_fifo_sink_eop;
wire [255:0] monroe_ionphoton_rtio_analyzer_fifo_sink_payload_data;
wire monroe_ionphoton_rtio_analyzer_fifo_source_stb;
wire monroe_ionphoton_rtio_analyzer_fifo_source_ack;
wire monroe_ionphoton_rtio_analyzer_fifo_source_eop;
wire [255:0] monroe_ionphoton_rtio_analyzer_fifo_source_payload_data;
wire monroe_ionphoton_rtio_analyzer_fifo_re;
reg monroe_ionphoton_rtio_analyzer_fifo_readable = 1'd0;
wire monroe_ionphoton_rtio_analyzer_fifo_syncfifo_we;
wire monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable;
wire monroe_ionphoton_rtio_analyzer_fifo_syncfifo_re;
wire monroe_ionphoton_rtio_analyzer_fifo_syncfifo_readable;
wire [256:0] monroe_ionphoton_rtio_analyzer_fifo_syncfifo_din;
wire [256:0] monroe_ionphoton_rtio_analyzer_fifo_syncfifo_dout;
reg [7:0] monroe_ionphoton_rtio_analyzer_fifo_level0 = 8'd0;
reg monroe_ionphoton_rtio_analyzer_fifo_replace = 1'd0;
reg [6:0] monroe_ionphoton_rtio_analyzer_fifo_produce = 7'd0;
reg [6:0] monroe_ionphoton_rtio_analyzer_fifo_consume = 7'd0;
reg [6:0] monroe_ionphoton_rtio_analyzer_fifo_wrport_adr;
wire [256:0] monroe_ionphoton_rtio_analyzer_fifo_wrport_dat_r;
wire monroe_ionphoton_rtio_analyzer_fifo_wrport_we;
wire [256:0] monroe_ionphoton_rtio_analyzer_fifo_wrport_dat_w;
wire monroe_ionphoton_rtio_analyzer_fifo_do_read;
wire [6:0] monroe_ionphoton_rtio_analyzer_fifo_rdport_adr;
wire [256:0] monroe_ionphoton_rtio_analyzer_fifo_rdport_dat_r;
wire monroe_ionphoton_rtio_analyzer_fifo_rdport_re;
wire [7:0] monroe_ionphoton_rtio_analyzer_fifo_level1;
wire [255:0] monroe_ionphoton_rtio_analyzer_fifo_fifo_in_payload_data;
wire monroe_ionphoton_rtio_analyzer_fifo_fifo_in_eop;
wire [255:0] monroe_ionphoton_rtio_analyzer_fifo_fifo_out_payload_data;
wire monroe_ionphoton_rtio_analyzer_fifo_fifo_out_eop;
wire monroe_ionphoton_rtio_analyzer_converter_sink_stb;
wire monroe_ionphoton_rtio_analyzer_converter_sink_ack;
wire monroe_ionphoton_rtio_analyzer_converter_sink_eop;
wire [255:0] monroe_ionphoton_rtio_analyzer_converter_sink_payload_data;
wire monroe_ionphoton_rtio_analyzer_converter_source_stb;
wire monroe_ionphoton_rtio_analyzer_converter_source_ack;
wire monroe_ionphoton_rtio_analyzer_converter_source_eop;
reg [127:0] monroe_ionphoton_rtio_analyzer_converter_source_payload_data;
wire monroe_ionphoton_rtio_analyzer_converter_source_payload_valid_token_count;
reg monroe_ionphoton_rtio_analyzer_converter_mux = 1'd0;
wire monroe_ionphoton_rtio_analyzer_converter_last;
wire monroe_ionphoton_rtio_analyzer_dma_reset_re;
wire monroe_ionphoton_rtio_analyzer_dma_reset_r;
reg monroe_ionphoton_rtio_analyzer_dma_reset_w = 1'd0;
reg [33:0] monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full = 34'd0;
wire [29:0] monroe_ionphoton_rtio_analyzer_dma_base_address_storage;
reg monroe_ionphoton_rtio_analyzer_dma_base_address_re = 1'd0;
reg [33:0] monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full = 34'd0;
wire [29:0] monroe_ionphoton_rtio_analyzer_dma_last_address_storage;
reg monroe_ionphoton_rtio_analyzer_dma_last_address_re = 1'd0;
wire [63:0] monroe_ionphoton_rtio_analyzer_dma_status;
wire monroe_ionphoton_rtio_analyzer_dma_sink_stb;
wire monroe_ionphoton_rtio_analyzer_dma_sink_ack;
wire monroe_ionphoton_rtio_analyzer_dma_sink_eop;
wire [127:0] monroe_ionphoton_rtio_analyzer_dma_sink_payload_data;
wire monroe_ionphoton_rtio_analyzer_dma_sink_payload_valid_token_count;
reg [58:0] monroe_ionphoton_rtio_analyzer_dma_message_count = 59'd0;
reg monroe_ionphoton_rtio_analyzer_enable_r = 1'd0;
reg [5:0] minicon_state = 6'd0;
reg [5:0] minicon_next_state;
reg [2:0] fullmemorywe_state = 3'd0;
reg [2:0] fullmemorywe_next_state;
reg [2:0] a7_1000basex_transmitpath_state = 3'd0;
reg [2:0] a7_1000basex_transmitpath_next_state;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value;
reg monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value_ce;
reg [2:0] a7_1000basex_receivepath_state = 3'd0;
reg [2:0] a7_1000basex_receivepath_next_state;
reg [1:0] a7_1000basex_fsm_state = 2'd0;
reg [1:0] a7_1000basex_fsm_next_state;
reg [1:0] a7_1000basex_gtptxinit_state = 2'd0;
reg [1:0] a7_1000basex_gtptxinit_next_state;
reg [3:0] a7_1000basex_gtprxinit_state = 4'd0;
reg [3:0] a7_1000basex_gtprxinit_next_state;
reg [15:0] monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value;
reg monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value_ce;
reg liteethmacgap_state = 1'd0;
reg liteethmacgap_next_state;
reg [1:0] liteethmacpreambleinserter_state = 2'd0;
reg [1:0] liteethmacpreambleinserter_next_state;
reg liteethmacpreamblechecker_state = 1'd0;
reg liteethmacpreamblechecker_next_state;
reg [1:0] liteethmaccrc32inserter_state = 2'd0;
reg [1:0] liteethmaccrc32inserter_next_state;
reg [1:0] liteethmaccrc32checker_state = 2'd0;
reg [1:0] liteethmaccrc32checker_next_state;
reg liteethmacpaddinginserter_state = 1'd0;
reg liteethmacpaddinginserter_next_state;
reg [1:0] liteethmacsramwriter_state = 2'd0;
reg [1:0] liteethmacsramwriter_next_state;
reg [31:0] monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value;
reg monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value_ce;
reg [1:0] liteethmacsramreader_state = 2'd0;
reg [1:0] liteethmacsramreader_next_state;
wire [29:0] shared_adr;
wire [31:0] shared_dat_w;
wire [31:0] shared_dat_r;
wire [3:0] shared_sel;
wire shared_cyc;
wire shared_stb;
wire shared_ack;
wire shared_we;
wire [2:0] shared_cti;
wire [1:0] shared_bte;
wire shared_err;
wire [1:0] request;
reg grant = 1'd0;
reg [4:0] slave_sel;
reg [4:0] slave_sel_r = 5'd0;
reg [2:0] spimaster0_state = 3'd0;
reg [2:0] spimaster0_next_state;
reg [2:0] spimaster1_state = 3'd0;
reg [2:0] spimaster1_next_state;
reg [2:0] spimaster2_state = 3'd0;
reg [2:0] spimaster2_next_state;
reg [1:0] clockdomainsrenamer_resetinserter_state = 2'd0;
reg [1:0] clockdomainsrenamer_resetinserter_next_state;
reg [1:0] clockdomainsrenamer_recordconverter_state = 2'd0;
reg [1:0] clockdomainsrenamer_recordconverter_next_state;
reg [2:0] clockdomainsrenamer_crimaster_state = 3'd0;
reg [2:0] clockdomainsrenamer_crimaster_next_state;
reg [2:0] clockdomainsrenamer_fsm_state = 3'd0;
reg [2:0] clockdomainsrenamer_fsm_next_state;
wire [1:0] sdram_cpulevel_arbiter_request;
reg sdram_cpulevel_arbiter_grant = 1'd0;
wire [2:0] sdram_native_arbiter_request;
reg [1:0] sdram_native_arbiter_grant = 2'd0;
wire [29:0] monroe_ionphoton_shared_adr;
wire [31:0] monroe_ionphoton_shared_dat_w;
wire [31:0] monroe_ionphoton_shared_dat_r;
wire [3:0] monroe_ionphoton_shared_sel;
wire monroe_ionphoton_shared_cyc;
wire monroe_ionphoton_shared_stb;
wire monroe_ionphoton_shared_ack;
wire monroe_ionphoton_shared_we;
wire [2:0] monroe_ionphoton_shared_cti;
wire [1:0] monroe_ionphoton_shared_bte;
wire monroe_ionphoton_shared_err;
wire [1:0] monroe_ionphoton_request;
reg monroe_ionphoton_grant = 1'd0;
reg [5:0] monroe_ionphoton_slave_sel;
reg [5:0] monroe_ionphoton_slave_sel_r = 6'd0;
wire [13:0] monroe_ionphoton_interface0_bank_bus_adr;
wire monroe_ionphoton_interface0_bank_bus_we;
wire [7:0] monroe_ionphoton_interface0_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface0_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank0_dly_sel0_re;
wire [1:0] monroe_ionphoton_csrbank0_dly_sel0_r;
wire [1:0] monroe_ionphoton_csrbank0_dly_sel0_w;
wire monroe_ionphoton_csrbank0_sel;
wire [13:0] monroe_ionphoton_interface1_bank_bus_adr;
wire monroe_ionphoton_interface1_bank_bus_we;
wire [7:0] monroe_ionphoton_interface1_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface1_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank1_control0_re;
wire [3:0] monroe_ionphoton_csrbank1_control0_r;
wire [3:0] monroe_ionphoton_csrbank1_control0_w;
wire monroe_ionphoton_csrbank1_pi0_command0_re;
wire [5:0] monroe_ionphoton_csrbank1_pi0_command0_r;
wire [5:0] monroe_ionphoton_csrbank1_pi0_command0_w;
wire monroe_ionphoton_csrbank1_pi0_address1_re;
wire [6:0] monroe_ionphoton_csrbank1_pi0_address1_r;
wire [6:0] monroe_ionphoton_csrbank1_pi0_address1_w;
wire monroe_ionphoton_csrbank1_pi0_address0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_address0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_address0_w;
wire monroe_ionphoton_csrbank1_pi0_baddress0_re;
wire [2:0] monroe_ionphoton_csrbank1_pi0_baddress0_r;
wire [2:0] monroe_ionphoton_csrbank1_pi0_baddress0_w;
wire monroe_ionphoton_csrbank1_pi0_wrdata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata3_w;
wire monroe_ionphoton_csrbank1_pi0_wrdata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata2_w;
wire monroe_ionphoton_csrbank1_pi0_wrdata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata1_w;
wire monroe_ionphoton_csrbank1_pi0_wrdata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_wrdata0_w;
wire monroe_ionphoton_csrbank1_pi0_rddata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata3_w;
wire monroe_ionphoton_csrbank1_pi0_rddata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata2_w;
wire monroe_ionphoton_csrbank1_pi0_rddata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata1_w;
wire monroe_ionphoton_csrbank1_pi0_rddata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi0_rddata0_w;
wire monroe_ionphoton_csrbank1_pi1_command0_re;
wire [5:0] monroe_ionphoton_csrbank1_pi1_command0_r;
wire [5:0] monroe_ionphoton_csrbank1_pi1_command0_w;
wire monroe_ionphoton_csrbank1_pi1_address1_re;
wire [6:0] monroe_ionphoton_csrbank1_pi1_address1_r;
wire [6:0] monroe_ionphoton_csrbank1_pi1_address1_w;
wire monroe_ionphoton_csrbank1_pi1_address0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_address0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_address0_w;
wire monroe_ionphoton_csrbank1_pi1_baddress0_re;
wire [2:0] monroe_ionphoton_csrbank1_pi1_baddress0_r;
wire [2:0] monroe_ionphoton_csrbank1_pi1_baddress0_w;
wire monroe_ionphoton_csrbank1_pi1_wrdata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata3_w;
wire monroe_ionphoton_csrbank1_pi1_wrdata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata2_w;
wire monroe_ionphoton_csrbank1_pi1_wrdata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata1_w;
wire monroe_ionphoton_csrbank1_pi1_wrdata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_wrdata0_w;
wire monroe_ionphoton_csrbank1_pi1_rddata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata3_w;
wire monroe_ionphoton_csrbank1_pi1_rddata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata2_w;
wire monroe_ionphoton_csrbank1_pi1_rddata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata1_w;
wire monroe_ionphoton_csrbank1_pi1_rddata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi1_rddata0_w;
wire monroe_ionphoton_csrbank1_pi2_command0_re;
wire [5:0] monroe_ionphoton_csrbank1_pi2_command0_r;
wire [5:0] monroe_ionphoton_csrbank1_pi2_command0_w;
wire monroe_ionphoton_csrbank1_pi2_address1_re;
wire [6:0] monroe_ionphoton_csrbank1_pi2_address1_r;
wire [6:0] monroe_ionphoton_csrbank1_pi2_address1_w;
wire monroe_ionphoton_csrbank1_pi2_address0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_address0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_address0_w;
wire monroe_ionphoton_csrbank1_pi2_baddress0_re;
wire [2:0] monroe_ionphoton_csrbank1_pi2_baddress0_r;
wire [2:0] monroe_ionphoton_csrbank1_pi2_baddress0_w;
wire monroe_ionphoton_csrbank1_pi2_wrdata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata3_w;
wire monroe_ionphoton_csrbank1_pi2_wrdata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata2_w;
wire monroe_ionphoton_csrbank1_pi2_wrdata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata1_w;
wire monroe_ionphoton_csrbank1_pi2_wrdata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_wrdata0_w;
wire monroe_ionphoton_csrbank1_pi2_rddata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata3_w;
wire monroe_ionphoton_csrbank1_pi2_rddata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata2_w;
wire monroe_ionphoton_csrbank1_pi2_rddata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata1_w;
wire monroe_ionphoton_csrbank1_pi2_rddata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi2_rddata0_w;
wire monroe_ionphoton_csrbank1_pi3_command0_re;
wire [5:0] monroe_ionphoton_csrbank1_pi3_command0_r;
wire [5:0] monroe_ionphoton_csrbank1_pi3_command0_w;
wire monroe_ionphoton_csrbank1_pi3_address1_re;
wire [6:0] monroe_ionphoton_csrbank1_pi3_address1_r;
wire [6:0] monroe_ionphoton_csrbank1_pi3_address1_w;
wire monroe_ionphoton_csrbank1_pi3_address0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_address0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_address0_w;
wire monroe_ionphoton_csrbank1_pi3_baddress0_re;
wire [2:0] monroe_ionphoton_csrbank1_pi3_baddress0_r;
wire [2:0] monroe_ionphoton_csrbank1_pi3_baddress0_w;
wire monroe_ionphoton_csrbank1_pi3_wrdata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata3_w;
wire monroe_ionphoton_csrbank1_pi3_wrdata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata2_w;
wire monroe_ionphoton_csrbank1_pi3_wrdata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata1_w;
wire monroe_ionphoton_csrbank1_pi3_wrdata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_wrdata0_w;
wire monroe_ionphoton_csrbank1_pi3_rddata3_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata3_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata3_w;
wire monroe_ionphoton_csrbank1_pi3_rddata2_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata2_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata2_w;
wire monroe_ionphoton_csrbank1_pi3_rddata1_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata1_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata1_w;
wire monroe_ionphoton_csrbank1_pi3_rddata0_re;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata0_r;
wire [7:0] monroe_ionphoton_csrbank1_pi3_rddata0_w;
wire monroe_ionphoton_csrbank1_sel;
wire [13:0] monroe_ionphoton_interface2_bank_bus_adr;
wire monroe_ionphoton_interface2_bank_bus_we;
wire [7:0] monroe_ionphoton_interface2_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface2_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank2_sram_writer_slot_re;
wire [1:0] monroe_ionphoton_csrbank2_sram_writer_slot_r;
wire [1:0] monroe_ionphoton_csrbank2_sram_writer_slot_w;
wire monroe_ionphoton_csrbank2_sram_writer_length3_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length3_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length3_w;
wire monroe_ionphoton_csrbank2_sram_writer_length2_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length2_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length2_w;
wire monroe_ionphoton_csrbank2_sram_writer_length1_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length1_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length1_w;
wire monroe_ionphoton_csrbank2_sram_writer_length0_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length0_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_length0_w;
wire monroe_ionphoton_csrbank2_sram_writer_errors3_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors3_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors3_w;
wire monroe_ionphoton_csrbank2_sram_writer_errors2_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors2_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors2_w;
wire monroe_ionphoton_csrbank2_sram_writer_errors1_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors1_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors1_w;
wire monroe_ionphoton_csrbank2_sram_writer_errors0_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors0_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_writer_errors0_w;
wire monroe_ionphoton_csrbank2_sram_writer_ev_enable0_re;
wire monroe_ionphoton_csrbank2_sram_writer_ev_enable0_r;
wire monroe_ionphoton_csrbank2_sram_writer_ev_enable0_w;
wire monroe_ionphoton_csrbank2_sram_reader_ready_re;
wire monroe_ionphoton_csrbank2_sram_reader_ready_r;
wire monroe_ionphoton_csrbank2_sram_reader_ready_w;
wire monroe_ionphoton_csrbank2_sram_reader_slot0_re;
wire [1:0] monroe_ionphoton_csrbank2_sram_reader_slot0_r;
wire [1:0] monroe_ionphoton_csrbank2_sram_reader_slot0_w;
wire monroe_ionphoton_csrbank2_sram_reader_length1_re;
wire [2:0] monroe_ionphoton_csrbank2_sram_reader_length1_r;
wire [2:0] monroe_ionphoton_csrbank2_sram_reader_length1_w;
wire monroe_ionphoton_csrbank2_sram_reader_length0_re;
wire [7:0] monroe_ionphoton_csrbank2_sram_reader_length0_r;
wire [7:0] monroe_ionphoton_csrbank2_sram_reader_length0_w;
wire monroe_ionphoton_csrbank2_sram_reader_ev_enable0_re;
wire monroe_ionphoton_csrbank2_sram_reader_ev_enable0_r;
wire monroe_ionphoton_csrbank2_sram_reader_ev_enable0_w;
wire monroe_ionphoton_csrbank2_preamble_errors3_re;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors3_r;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors3_w;
wire monroe_ionphoton_csrbank2_preamble_errors2_re;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors2_r;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors2_w;
wire monroe_ionphoton_csrbank2_preamble_errors1_re;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors1_r;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors1_w;
wire monroe_ionphoton_csrbank2_preamble_errors0_re;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors0_r;
wire [7:0] monroe_ionphoton_csrbank2_preamble_errors0_w;
wire monroe_ionphoton_csrbank2_crc_errors3_re;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors3_r;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors3_w;
wire monroe_ionphoton_csrbank2_crc_errors2_re;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors2_r;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors2_w;
wire monroe_ionphoton_csrbank2_crc_errors1_re;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors1_r;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors1_w;
wire monroe_ionphoton_csrbank2_crc_errors0_re;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors0_r;
wire [7:0] monroe_ionphoton_csrbank2_crc_errors0_w;
wire monroe_ionphoton_csrbank2_sel;
wire [13:0] monroe_ionphoton_interface3_bank_bus_adr;
wire monroe_ionphoton_interface3_bank_bus_we;
wire [7:0] monroe_ionphoton_interface3_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface3_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank3_in_re;
wire [1:0] monroe_ionphoton_csrbank3_in_r;
wire [1:0] monroe_ionphoton_csrbank3_in_w;
wire monroe_ionphoton_csrbank3_out0_re;
wire [1:0] monroe_ionphoton_csrbank3_out0_r;
wire [1:0] monroe_ionphoton_csrbank3_out0_w;
wire monroe_ionphoton_csrbank3_oe0_re;
wire [1:0] monroe_ionphoton_csrbank3_oe0_r;
wire [1:0] monroe_ionphoton_csrbank3_oe0_w;
wire monroe_ionphoton_csrbank3_sel;
wire [13:0] monroe_ionphoton_interface4_bank_bus_adr;
wire monroe_ionphoton_interface4_bank_bus_we;
wire [7:0] monroe_ionphoton_interface4_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface4_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank4_address0_re;
wire [7:0] monroe_ionphoton_csrbank4_address0_r;
wire [7:0] monroe_ionphoton_csrbank4_address0_w;
wire monroe_ionphoton_csrbank4_data_re;
wire [7:0] monroe_ionphoton_csrbank4_data_r;
wire [7:0] monroe_ionphoton_csrbank4_data_w;
wire monroe_ionphoton_csrbank4_sel;
wire [13:0] monroe_ionphoton_interface5_bank_bus_adr;
wire monroe_ionphoton_interface5_bank_bus_we;
wire [7:0] monroe_ionphoton_interface5_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface5_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank5_reset0_re;
wire monroe_ionphoton_csrbank5_reset0_r;
wire monroe_ionphoton_csrbank5_reset0_w;
wire monroe_ionphoton_csrbank5_sel;
wire [13:0] monroe_ionphoton_interface6_bank_bus_adr;
wire monroe_ionphoton_interface6_bank_bus_we;
wire [7:0] monroe_ionphoton_interface6_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface6_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank6_out0_re;
wire monroe_ionphoton_csrbank6_out0_r;
wire monroe_ionphoton_csrbank6_out0_w;
wire monroe_ionphoton_csrbank6_sel;
wire [13:0] monroe_ionphoton_interface7_bank_bus_adr;
wire monroe_ionphoton_interface7_bank_bus_we;
wire [7:0] monroe_ionphoton_interface7_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface7_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank7_enable0_re;
wire monroe_ionphoton_csrbank7_enable0_r;
wire monroe_ionphoton_csrbank7_enable0_w;
wire monroe_ionphoton_csrbank7_busy_re;
wire monroe_ionphoton_csrbank7_busy_r;
wire monroe_ionphoton_csrbank7_busy_w;
wire monroe_ionphoton_csrbank7_message_encoder_overflow_re;
wire monroe_ionphoton_csrbank7_message_encoder_overflow_r;
wire monroe_ionphoton_csrbank7_message_encoder_overflow_w;
wire monroe_ionphoton_csrbank7_dma_base_address4_re;
wire [1:0] monroe_ionphoton_csrbank7_dma_base_address4_r;
wire [1:0] monroe_ionphoton_csrbank7_dma_base_address4_w;
wire monroe_ionphoton_csrbank7_dma_base_address3_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address3_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address3_w;
wire monroe_ionphoton_csrbank7_dma_base_address2_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address2_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address2_w;
wire monroe_ionphoton_csrbank7_dma_base_address1_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address1_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address1_w;
wire monroe_ionphoton_csrbank7_dma_base_address0_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address0_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_base_address0_w;
wire monroe_ionphoton_csrbank7_dma_last_address4_re;
wire [1:0] monroe_ionphoton_csrbank7_dma_last_address4_r;
wire [1:0] monroe_ionphoton_csrbank7_dma_last_address4_w;
wire monroe_ionphoton_csrbank7_dma_last_address3_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address3_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address3_w;
wire monroe_ionphoton_csrbank7_dma_last_address2_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address2_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address2_w;
wire monroe_ionphoton_csrbank7_dma_last_address1_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address1_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address1_w;
wire monroe_ionphoton_csrbank7_dma_last_address0_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address0_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_last_address0_w;
wire monroe_ionphoton_csrbank7_dma_byte_count7_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count7_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count7_w;
wire monroe_ionphoton_csrbank7_dma_byte_count6_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count6_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count6_w;
wire monroe_ionphoton_csrbank7_dma_byte_count5_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count5_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count5_w;
wire monroe_ionphoton_csrbank7_dma_byte_count4_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count4_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count4_w;
wire monroe_ionphoton_csrbank7_dma_byte_count3_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count3_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count3_w;
wire monroe_ionphoton_csrbank7_dma_byte_count2_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count2_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count2_w;
wire monroe_ionphoton_csrbank7_dma_byte_count1_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count1_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count1_w;
wire monroe_ionphoton_csrbank7_dma_byte_count0_re;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count0_r;
wire [7:0] monroe_ionphoton_csrbank7_dma_byte_count0_w;
wire monroe_ionphoton_csrbank7_sel;
wire [13:0] monroe_ionphoton_interface8_bank_bus_adr;
wire monroe_ionphoton_interface8_bank_bus_we;
wire [7:0] monroe_ionphoton_interface8_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface8_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank8_collision_channel1_re;
wire [7:0] monroe_ionphoton_csrbank8_collision_channel1_r;
wire [7:0] monroe_ionphoton_csrbank8_collision_channel1_w;
wire monroe_ionphoton_csrbank8_collision_channel0_re;
wire [7:0] monroe_ionphoton_csrbank8_collision_channel0_r;
wire [7:0] monroe_ionphoton_csrbank8_collision_channel0_w;
wire monroe_ionphoton_csrbank8_busy_channel1_re;
wire [7:0] monroe_ionphoton_csrbank8_busy_channel1_r;
wire [7:0] monroe_ionphoton_csrbank8_busy_channel1_w;
wire monroe_ionphoton_csrbank8_busy_channel0_re;
wire [7:0] monroe_ionphoton_csrbank8_busy_channel0_r;
wire [7:0] monroe_ionphoton_csrbank8_busy_channel0_w;
wire monroe_ionphoton_csrbank8_sequence_error_channel1_re;
wire [7:0] monroe_ionphoton_csrbank8_sequence_error_channel1_r;
wire [7:0] monroe_ionphoton_csrbank8_sequence_error_channel1_w;
wire monroe_ionphoton_csrbank8_sequence_error_channel0_re;
wire [7:0] monroe_ionphoton_csrbank8_sequence_error_channel0_r;
wire [7:0] monroe_ionphoton_csrbank8_sequence_error_channel0_w;
wire monroe_ionphoton_csrbank8_sel;
wire [13:0] monroe_ionphoton_interface9_bank_bus_adr;
wire monroe_ionphoton_interface9_bank_bus_we;
wire [7:0] monroe_ionphoton_interface9_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface9_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank9_pll_reset0_re;
wire monroe_ionphoton_csrbank9_pll_reset0_r;
wire monroe_ionphoton_csrbank9_pll_reset0_w;
wire monroe_ionphoton_csrbank9_pll_locked_re;
wire monroe_ionphoton_csrbank9_pll_locked_r;
wire monroe_ionphoton_csrbank9_pll_locked_w;
wire monroe_ionphoton_csrbank9_sel;
wire [13:0] monroe_ionphoton_interface10_bank_bus_adr;
wire monroe_ionphoton_interface10_bank_bus_we;
wire [7:0] monroe_ionphoton_interface10_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface10_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank10_mon_chan_sel0_re;
wire [5:0] monroe_ionphoton_csrbank10_mon_chan_sel0_r;
wire [5:0] monroe_ionphoton_csrbank10_mon_chan_sel0_w;
wire monroe_ionphoton_csrbank10_mon_probe_sel0_re;
wire monroe_ionphoton_csrbank10_mon_probe_sel0_r;
wire monroe_ionphoton_csrbank10_mon_probe_sel0_w;
wire monroe_ionphoton_csrbank10_mon_value_re;
wire monroe_ionphoton_csrbank10_mon_value_r;
wire monroe_ionphoton_csrbank10_mon_value_w;
wire monroe_ionphoton_csrbank10_inj_chan_sel0_re;
wire [5:0] monroe_ionphoton_csrbank10_inj_chan_sel0_r;
wire [5:0] monroe_ionphoton_csrbank10_inj_chan_sel0_w;
wire monroe_ionphoton_csrbank10_inj_override_sel0_re;
wire [1:0] monroe_ionphoton_csrbank10_inj_override_sel0_r;
wire [1:0] monroe_ionphoton_csrbank10_inj_override_sel0_w;
wire monroe_ionphoton_csrbank10_sel;
wire [13:0] monroe_ionphoton_interface11_bank_bus_adr;
wire monroe_ionphoton_interface11_bank_bus_we;
wire [7:0] monroe_ionphoton_interface11_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface11_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank11_bitbang0_re;
wire [3:0] monroe_ionphoton_csrbank11_bitbang0_r;
wire [3:0] monroe_ionphoton_csrbank11_bitbang0_w;
wire monroe_ionphoton_csrbank11_miso_re;
wire monroe_ionphoton_csrbank11_miso_r;
wire monroe_ionphoton_csrbank11_miso_w;
wire monroe_ionphoton_csrbank11_bitbang_en0_re;
wire monroe_ionphoton_csrbank11_bitbang_en0_r;
wire monroe_ionphoton_csrbank11_bitbang_en0_w;
wire monroe_ionphoton_csrbank11_sel;
wire [13:0] monroe_ionphoton_interface12_bank_bus_adr;
wire monroe_ionphoton_interface12_bank_bus_we;
wire [7:0] monroe_ionphoton_interface12_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface12_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank12_load7_re;
wire [7:0] monroe_ionphoton_csrbank12_load7_r;
wire [7:0] monroe_ionphoton_csrbank12_load7_w;
wire monroe_ionphoton_csrbank12_load6_re;
wire [7:0] monroe_ionphoton_csrbank12_load6_r;
wire [7:0] monroe_ionphoton_csrbank12_load6_w;
wire monroe_ionphoton_csrbank12_load5_re;
wire [7:0] monroe_ionphoton_csrbank12_load5_r;
wire [7:0] monroe_ionphoton_csrbank12_load5_w;
wire monroe_ionphoton_csrbank12_load4_re;
wire [7:0] monroe_ionphoton_csrbank12_load4_r;
wire [7:0] monroe_ionphoton_csrbank12_load4_w;
wire monroe_ionphoton_csrbank12_load3_re;
wire [7:0] monroe_ionphoton_csrbank12_load3_r;
wire [7:0] monroe_ionphoton_csrbank12_load3_w;
wire monroe_ionphoton_csrbank12_load2_re;
wire [7:0] monroe_ionphoton_csrbank12_load2_r;
wire [7:0] monroe_ionphoton_csrbank12_load2_w;
wire monroe_ionphoton_csrbank12_load1_re;
wire [7:0] monroe_ionphoton_csrbank12_load1_r;
wire [7:0] monroe_ionphoton_csrbank12_load1_w;
wire monroe_ionphoton_csrbank12_load0_re;
wire [7:0] monroe_ionphoton_csrbank12_load0_r;
wire [7:0] monroe_ionphoton_csrbank12_load0_w;
wire monroe_ionphoton_csrbank12_reload7_re;
wire [7:0] monroe_ionphoton_csrbank12_reload7_r;
wire [7:0] monroe_ionphoton_csrbank12_reload7_w;
wire monroe_ionphoton_csrbank12_reload6_re;
wire [7:0] monroe_ionphoton_csrbank12_reload6_r;
wire [7:0] monroe_ionphoton_csrbank12_reload6_w;
wire monroe_ionphoton_csrbank12_reload5_re;
wire [7:0] monroe_ionphoton_csrbank12_reload5_r;
wire [7:0] monroe_ionphoton_csrbank12_reload5_w;
wire monroe_ionphoton_csrbank12_reload4_re;
wire [7:0] monroe_ionphoton_csrbank12_reload4_r;
wire [7:0] monroe_ionphoton_csrbank12_reload4_w;
wire monroe_ionphoton_csrbank12_reload3_re;
wire [7:0] monroe_ionphoton_csrbank12_reload3_r;
wire [7:0] monroe_ionphoton_csrbank12_reload3_w;
wire monroe_ionphoton_csrbank12_reload2_re;
wire [7:0] monroe_ionphoton_csrbank12_reload2_r;
wire [7:0] monroe_ionphoton_csrbank12_reload2_w;
wire monroe_ionphoton_csrbank12_reload1_re;
wire [7:0] monroe_ionphoton_csrbank12_reload1_r;
wire [7:0] monroe_ionphoton_csrbank12_reload1_w;
wire monroe_ionphoton_csrbank12_reload0_re;
wire [7:0] monroe_ionphoton_csrbank12_reload0_r;
wire [7:0] monroe_ionphoton_csrbank12_reload0_w;
wire monroe_ionphoton_csrbank12_en0_re;
wire monroe_ionphoton_csrbank12_en0_r;
wire monroe_ionphoton_csrbank12_en0_w;
wire monroe_ionphoton_csrbank12_value7_re;
wire [7:0] monroe_ionphoton_csrbank12_value7_r;
wire [7:0] monroe_ionphoton_csrbank12_value7_w;
wire monroe_ionphoton_csrbank12_value6_re;
wire [7:0] monroe_ionphoton_csrbank12_value6_r;
wire [7:0] monroe_ionphoton_csrbank12_value6_w;
wire monroe_ionphoton_csrbank12_value5_re;
wire [7:0] monroe_ionphoton_csrbank12_value5_r;
wire [7:0] monroe_ionphoton_csrbank12_value5_w;
wire monroe_ionphoton_csrbank12_value4_re;
wire [7:0] monroe_ionphoton_csrbank12_value4_r;
wire [7:0] monroe_ionphoton_csrbank12_value4_w;
wire monroe_ionphoton_csrbank12_value3_re;
wire [7:0] monroe_ionphoton_csrbank12_value3_r;
wire [7:0] monroe_ionphoton_csrbank12_value3_w;
wire monroe_ionphoton_csrbank12_value2_re;
wire [7:0] monroe_ionphoton_csrbank12_value2_r;
wire [7:0] monroe_ionphoton_csrbank12_value2_w;
wire monroe_ionphoton_csrbank12_value1_re;
wire [7:0] monroe_ionphoton_csrbank12_value1_r;
wire [7:0] monroe_ionphoton_csrbank12_value1_w;
wire monroe_ionphoton_csrbank12_value0_re;
wire [7:0] monroe_ionphoton_csrbank12_value0_r;
wire [7:0] monroe_ionphoton_csrbank12_value0_w;
wire monroe_ionphoton_csrbank12_ev_enable0_re;
wire monroe_ionphoton_csrbank12_ev_enable0_r;
wire monroe_ionphoton_csrbank12_ev_enable0_w;
wire monroe_ionphoton_csrbank12_sel;
wire [13:0] monroe_ionphoton_interface13_bank_bus_adr;
wire monroe_ionphoton_interface13_bank_bus_we;
wire [7:0] monroe_ionphoton_interface13_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface13_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank13_enable_null0_re;
wire monroe_ionphoton_csrbank13_enable_null0_r;
wire monroe_ionphoton_csrbank13_enable_null0_w;
wire monroe_ionphoton_csrbank13_enable_prog0_re;
wire monroe_ionphoton_csrbank13_enable_prog0_r;
wire monroe_ionphoton_csrbank13_enable_prog0_w;
wire monroe_ionphoton_csrbank13_prog_address3_re;
wire [5:0] monroe_ionphoton_csrbank13_prog_address3_r;
wire [5:0] monroe_ionphoton_csrbank13_prog_address3_w;
wire monroe_ionphoton_csrbank13_prog_address2_re;
wire [7:0] monroe_ionphoton_csrbank13_prog_address2_r;
wire [7:0] monroe_ionphoton_csrbank13_prog_address2_w;
wire monroe_ionphoton_csrbank13_prog_address1_re;
wire [7:0] monroe_ionphoton_csrbank13_prog_address1_r;
wire [7:0] monroe_ionphoton_csrbank13_prog_address1_w;
wire monroe_ionphoton_csrbank13_prog_address0_re;
wire [7:0] monroe_ionphoton_csrbank13_prog_address0_r;
wire [7:0] monroe_ionphoton_csrbank13_prog_address0_w;
wire monroe_ionphoton_csrbank13_sel;
wire [13:0] monroe_ionphoton_interface14_bank_bus_adr;
wire monroe_ionphoton_interface14_bank_bus_we;
wire [7:0] monroe_ionphoton_interface14_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface14_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank14_txfull_re;
wire monroe_ionphoton_csrbank14_txfull_r;
wire monroe_ionphoton_csrbank14_txfull_w;
wire monroe_ionphoton_csrbank14_rxempty_re;
wire monroe_ionphoton_csrbank14_rxempty_r;
wire monroe_ionphoton_csrbank14_rxempty_w;
wire monroe_ionphoton_csrbank14_ev_enable0_re;
wire [1:0] monroe_ionphoton_csrbank14_ev_enable0_r;
wire [1:0] monroe_ionphoton_csrbank14_ev_enable0_w;
wire monroe_ionphoton_csrbank14_sel;
wire [13:0] monroe_ionphoton_interface15_bank_bus_adr;
wire monroe_ionphoton_interface15_bank_bus_we;
wire [7:0] monroe_ionphoton_interface15_bank_bus_dat_w;
reg [7:0] monroe_ionphoton_interface15_bank_bus_dat_r = 8'd0;
wire monroe_ionphoton_csrbank15_tuning_word3_re;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word3_r;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word3_w;
wire monroe_ionphoton_csrbank15_tuning_word2_re;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word2_r;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word2_w;
wire monroe_ionphoton_csrbank15_tuning_word1_re;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word1_r;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word1_w;
wire monroe_ionphoton_csrbank15_tuning_word0_re;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word0_r;
wire [7:0] monroe_ionphoton_csrbank15_tuning_word0_w;
wire monroe_ionphoton_csrbank15_sel;
reg [29:0] comb_rhs_array_muxed0;
reg [31:0] comb_rhs_array_muxed1;
reg [3:0] comb_rhs_array_muxed2;
reg comb_rhs_array_muxed3;
reg comb_rhs_array_muxed4;
reg comb_rhs_array_muxed5;
reg [2:0] comb_rhs_array_muxed6;
reg [1:0] comb_rhs_array_muxed7;
wire comb_lhs_array_muxed;
reg comb_rhs_array_muxed8;
reg [1:0] comb_rhs_array_muxed9;
reg [1:0] comb_rhs_array_muxed10;
reg [23:0] comb_rhs_array_muxed11;
reg [63:0] comb_rhs_array_muxed12;
reg [511:0] comb_rhs_array_muxed13;
reg [7:0] comb_rhs_array_muxed14;
reg [63:0] comb_rhs_array_muxed15;
reg comb_rhs_array_muxed16;
reg comb_rhs_array_muxed17;
reg comb_rhs_array_muxed18;
reg comb_rhs_array_muxed19;
reg comb_rhs_array_muxed20;
reg comb_rhs_array_muxed21;
reg comb_rhs_array_muxed22;
reg comb_rhs_array_muxed23;
reg comb_rhs_array_muxed24;
reg comb_rhs_array_muxed25;
reg comb_rhs_array_muxed26;
reg comb_rhs_array_muxed27;
reg comb_rhs_array_muxed28;
reg comb_rhs_array_muxed29;
reg comb_rhs_array_muxed30;
reg comb_rhs_array_muxed31;
reg comb_rhs_array_muxed32;
reg comb_rhs_array_muxed33;
reg comb_rhs_array_muxed34;
reg comb_rhs_array_muxed35;
reg comb_rhs_array_muxed36;
reg comb_rhs_array_muxed37;
reg comb_rhs_array_muxed38;
reg comb_rhs_array_muxed39;
reg comb_rhs_array_muxed40;
reg comb_rhs_array_muxed41;
reg comb_rhs_array_muxed42;
reg comb_rhs_array_muxed43;
reg comb_rhs_array_muxed44;
reg comb_rhs_array_muxed45;
reg comb_rhs_array_muxed46;
reg comb_rhs_array_muxed47;
reg comb_rhs_array_muxed48;
reg comb_rhs_array_muxed49;
reg comb_rhs_array_muxed50;
reg comb_rhs_array_muxed51;
reg comb_rhs_array_muxed52;
reg comb_rhs_array_muxed53;
reg [29:0] comb_rhs_array_muxed54;
reg [31:0] comb_rhs_array_muxed55;
reg [3:0] comb_rhs_array_muxed56;
reg comb_rhs_array_muxed57;
reg comb_rhs_array_muxed58;
reg comb_rhs_array_muxed59;
reg [2:0] comb_rhs_array_muxed60;
reg [1:0] comb_rhs_array_muxed61;
reg [29:0] comb_rhs_array_muxed62;
reg [127:0] comb_rhs_array_muxed63;
reg [15:0] comb_rhs_array_muxed64;
reg comb_rhs_array_muxed65;
reg comb_rhs_array_muxed66;
reg comb_rhs_array_muxed67;
reg [2:0] comb_rhs_array_muxed68;
reg [1:0] comb_rhs_array_muxed69;
reg [29:0] comb_rhs_array_muxed70;
reg [31:0] comb_rhs_array_muxed71;
reg [3:0] comb_rhs_array_muxed72;
reg comb_rhs_array_muxed73;
reg comb_rhs_array_muxed74;
reg comb_rhs_array_muxed75;
reg [2:0] comb_rhs_array_muxed76;
reg [1:0] comb_rhs_array_muxed77;
reg [2:0] sync_t_rhs_array_muxed0;
reg [2:0] sync_f_t_array_muxed0;
reg [2:0] sync_f_rhs_array_muxed0;
reg [4:0] sync_rhs_array_muxed0;
reg [5:0] sync_f_rhs_array_muxed1;
reg sync_f_rhs_array_muxed2;
reg sync_f_rhs_array_muxed3;
reg [3:0] sync_rhs_array_muxed1;
reg sync_rhs_array_muxed2;
reg sync_f_rhs_array_muxed4;
reg sync_basiclowerer_array_muxed0;
reg sync_basiclowerer_array_muxed1;
reg sync_basiclowerer_array_muxed2;
reg sync_basiclowerer_array_muxed3;
reg sync_basiclowerer_array_muxed4;
reg sync_basiclowerer_array_muxed5;
reg sync_basiclowerer_array_muxed6;
reg sync_basiclowerer_array_muxed7;
reg [7:0] sync_f_t_array_muxed1;
reg [6:0] sync_f_t_array_muxed2;
reg [7:0] sync_f_t_array_muxed3;
reg [6:0] sync_f_t_array_muxed4;
reg [7:0] sync_f_t_array_muxed5;
reg [6:0] sync_f_t_array_muxed6;
reg [7:0] sync_f_t_array_muxed7;
reg [6:0] sync_f_t_array_muxed8;
reg [7:0] sync_f_t_array_muxed9;
reg [6:0] sync_f_t_array_muxed10;
reg [7:0] sync_f_t_array_muxed11;
reg [6:0] sync_f_t_array_muxed12;
reg [7:0] sync_f_t_array_muxed13;
reg [6:0] sync_f_t_array_muxed14;
reg [7:0] sync_f_t_array_muxed15;
reg [6:0] sync_f_t_array_muxed16;
reg [7:0] sync_f_t_array_muxed17;
reg [6:0] sync_f_t_array_muxed18;
reg [7:0] sync_f_t_array_muxed19;
reg [6:0] sync_f_t_array_muxed20;
reg [7:0] sync_f_t_array_muxed21;
reg [6:0] sync_f_t_array_muxed22;
reg [7:0] sync_f_t_array_muxed23;
reg [6:0] sync_f_t_array_muxed24;
reg [7:0] sync_f_t_array_muxed25;
reg [6:0] sync_f_t_array_muxed26;
reg [7:0] sync_f_t_array_muxed27;
reg [6:0] sync_f_t_array_muxed28;
reg [7:0] sync_f_t_array_muxed29;
reg [6:0] sync_f_t_array_muxed30;
reg [7:0] sync_f_t_array_muxed31;
reg [6:0] sync_f_t_array_muxed32;
reg [7:0] sync_f_t_array_muxed33;
reg [6:0] sync_f_t_array_muxed34;
reg [7:0] sync_f_t_array_muxed35;
reg [6:0] sync_f_t_array_muxed36;
reg [7:0] sync_f_t_array_muxed37;
reg [6:0] sync_f_t_array_muxed38;
reg [7:0] sync_f_t_array_muxed39;
reg [6:0] sync_f_t_array_muxed40;
reg [7:0] sync_f_t_array_muxed41;
reg [6:0] sync_f_t_array_muxed42;
reg [7:0] sync_f_t_array_muxed43;
reg [6:0] sync_f_t_array_muxed44;
reg [7:0] sync_f_t_array_muxed45;
reg [6:0] sync_f_t_array_muxed46;
reg [7:0] sync_f_t_array_muxed47;
reg [6:0] sync_f_t_array_muxed48;
reg [7:0] sync_f_t_array_muxed49;
reg [6:0] sync_f_t_array_muxed50;
reg [7:0] sync_f_t_array_muxed51;
reg [6:0] sync_f_t_array_muxed52;
reg [7:0] sync_f_t_array_muxed53;
reg [6:0] sync_f_t_array_muxed54;
reg [7:0] sync_f_t_array_muxed55;
reg [6:0] sync_f_t_array_muxed56;
reg [7:0] sync_f_t_array_muxed57;
reg [6:0] sync_f_t_array_muxed58;
reg [7:0] sync_f_t_array_muxed59;
reg [6:0] sync_f_t_array_muxed60;
reg [7:0] sync_f_t_array_muxed61;
reg [6:0] sync_f_t_array_muxed62;
reg [60:0] sync_rhs_array_muxed3;
reg [60:0] sync_rhs_array_muxed4;
reg [60:0] sync_t_lhs_array_muxed = 61'd0;
reg [31:0] sync_t_rhs_array_muxed1;
reg [64:0] sync_t_rhs_array_muxed2;
reg [31:0] sync_rhs_array_muxed5;
reg [31:0] sync_t_t_array_muxed0 = 32'd0;
reg [31:0] sync_rhs_array_muxed6;
reg [31:0] sync_t_t_array_muxed1 = 32'd0;
reg sync_t_rhs_array_muxed3;
reg sync_t_rhs_array_muxed4;
reg sync_t_rhs_array_muxed5;
reg sync_t_rhs_array_muxed6;
reg sync_t_rhs_array_muxed7;
reg sync_t_rhs_array_muxed8;
reg sync_t_rhs_array_muxed9;
reg sync_t_rhs_array_muxed10;
reg sync_t_rhs_array_muxed11;
reg sync_t_rhs_array_muxed12;
reg sync_t_rhs_array_muxed13;
reg sync_t_rhs_array_muxed14;
reg sync_t_rhs_array_muxed15;
reg sync_t_rhs_array_muxed16;
reg sync_t_rhs_array_muxed17;
reg sync_t_rhs_array_muxed18;
reg sync_t_rhs_array_muxed19;
reg sync_t_rhs_array_muxed20;
reg sync_t_rhs_array_muxed21;
reg sync_t_rhs_array_muxed22;
reg sync_t_rhs_array_muxed23;
reg sync_t_rhs_array_muxed24;
reg sync_t_rhs_array_muxed25;
reg sync_t_rhs_array_muxed26;
reg sync_t_rhs_array_muxed27;
reg sync_t_rhs_array_muxed28;
reg sync_t_rhs_array_muxed29;
reg sync_t_rhs_array_muxed30;
reg sync_t_rhs_array_muxed31;
reg sync_t_rhs_array_muxed32;
reg sync_t_rhs_array_muxed33;
reg sync_t_rhs_array_muxed34;
reg sync_t_rhs_array_muxed35;
reg sync_t_rhs_array_muxed36;
reg sync_t_rhs_array_muxed37;
reg sync_t_rhs_array_muxed38;
reg sync_t_rhs_array_muxed39;
reg sync_t_rhs_array_muxed40;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl0_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl0;
wire xilinxasyncresetsynchronizerimpl0_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl1_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl1_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl2_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl2_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl3_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl3_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl1;
wire xilinxasyncresetsynchronizerimpl1_rst_meta;
wire xilinxasyncresetsynchronizerimpl2;
wire xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl4_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl4_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl5_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl5_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl6_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl6_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl7_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl7_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl8_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl9_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl9_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl10_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl10_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl11_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl11_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl12_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl12_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl13_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl13_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl14_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl14_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl3;
wire xilinxasyncresetsynchronizerimpl3_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl15_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl15_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [60:0] xilinxmultiregimpl16_regs0 = 61'd0;
(* async_reg = "true", dont_touch = "true" *) reg [60:0] xilinxmultiregimpl16_regs1 = 61'd0;
wire xilinxasyncresetsynchronizerimpl4_rst_meta;
wire xilinxasyncresetsynchronizerimpl5_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl17_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl17_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl18_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl18_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl19_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl19_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl20_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl20_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl21_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl21_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl22_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl22_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl23_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl23_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl24_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl24_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl25_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl25_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl26_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl26_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl27_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl27_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl28_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl28_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl29_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl29_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl30_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl30_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl31_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl31_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl32_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] xilinxmultiregimpl32_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl33_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl33_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl34_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl34_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl36_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl36_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl37_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl37_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl38_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl38_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl39_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl39_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl40_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl40_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl41_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl41_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl42_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl42_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl43_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl43_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl44_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl44_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl45_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl45_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl46_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl46_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl47_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl47_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl48_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl48_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl49_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl49_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl50_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl50_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl51_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl51_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl52_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl52_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl53_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl53_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl54_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl54_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl55_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl55_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl56_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl56_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl57_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl57_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl58_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl58_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl59_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl59_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl60_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl60_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl61_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl61_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl62_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl62_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] xilinxmultiregimpl63_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] xilinxmultiregimpl63_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl64_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl64_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl65_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl65_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] xilinxmultiregimpl66_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] xilinxmultiregimpl66_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl67_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl67_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl68_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl68_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl69_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl69_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl70_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl70_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl71_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl71_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl72_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl72_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl73_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl73_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl74_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl74_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl75_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl75_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl76_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl76_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl77_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl77_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl78_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl78_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl79_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl79_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl80_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl80_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl81_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl81_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl82_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl82_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl83_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl83_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl84_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl84_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl85_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl85_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl86_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl86_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl87_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl87_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl88_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl88_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl89_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl89_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl90_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl90_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl91_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl91_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl92_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl92_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl93_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl93_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl94_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl94_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl95_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl95_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl96_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl96_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl97_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl97_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl98_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl98_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl99_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl99_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl100_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl100_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl101_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl101_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl102_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl102_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl103_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl103_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl104_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl104_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl105_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl105_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl106_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl106_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl107_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl107_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl108_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl108_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl109_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl109_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl110_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl110_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl111_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl111_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl112_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl112_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl113_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl113_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl114_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl114_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl115_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl115_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl116_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl116_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl117_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl117_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl118_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl118_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl119_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl119_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl120_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl120_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl121_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl121_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl122_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl122_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl123_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl123_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl124_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl124_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl125_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl125_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl126_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl126_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl127_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl127_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl128_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl128_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl129_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl129_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl130_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl130_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl131_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl131_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl132_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl132_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl133_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl133_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl134_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl134_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl135_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl135_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl136_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl136_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl137_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl137_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl138_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl138_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl139_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl139_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl140_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl140_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl141_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl141_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl142_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl142_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl143_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl143_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl144_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl144_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl145_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl145_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl146_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl146_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl147_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl147_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl148_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl148_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl149_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl149_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl150_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl150_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl151_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl151_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl152_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl152_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl153_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl153_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl154_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl154_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl155_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl155_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl156_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl156_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl157_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl157_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl158_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl158_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl159_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl159_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl160_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl160_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl161_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl161_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl162_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl162_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl163_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl163_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl164_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl164_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl165_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl165_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl166_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl166_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl167_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl167_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl168_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl168_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl169_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl169_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl170_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl170_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl171_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl171_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl172_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl172_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg xilinxmultiregimpl173_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl173_regs1 = 1'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_valid;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_bank;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cas_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cas_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cs_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cs_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_ras_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_ras_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_we_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_we_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cke;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_odt;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_reset_n;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_mask = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata_mask;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_en = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata_en;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata_valid = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_valid;
assign sfp_ctl_rate_select = 1'd0;
assign sfp_ctl_tx_disable = 1'd0;
assign sfp_ctl_led = ((((~sfp_ctl_los) & (~sfp_ctl_tx_fault)) & sfp_ctl_mod_present) & monroe_ionphoton_monroe_ionphoton_pcs_link_up);
assign clk_sel = 1'd1;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt[0] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_irq;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt[1] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_irq;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt[2] <= monroe_ionphoton_monroe_ionphoton_ev_irq;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_i_adr_o[31:2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_d_adr_o[31:2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_adr;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_sel = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_sel;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cyc = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cyc;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_we;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cti = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cti;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_bte = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_bte;

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_err <= 1'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_err <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_ack | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_err);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_ack <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_ack;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_err <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_err;
	end
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[0] <= (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel[0]);
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[1] <= (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel[1]);
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[2] <= (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel[2]);
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[3] <= (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel[3]);
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_adr[9:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_re;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_txfull_status = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_ack);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_ack = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_trigger = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_ack);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_ack = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxempty_status = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_stb);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_ack = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_clear;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_trigger = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_stb);

// synthesis translate_off
reg dummy_d_3;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_clear <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_r[0])) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_3 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_4;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_w <= 2'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_w[0] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_status;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_w[1] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_status;
// synthesis translate_off
	dummy_d_4 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_5;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_clear <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_r[1])) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_5 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_6;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w <= 2'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w[0] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_pending;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w[1] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_pending;
// synthesis translate_off
	dummy_d_6 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_irq = ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage[0]) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage[1]));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_status = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_trigger;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_status = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_trigger;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_din = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_payload_data};
assign {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_payload_data} = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_ack = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_in_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_fifo_out_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_re = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_7;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr <= 4'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_replace) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_7 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_we = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_we & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_replace));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_do_read = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_readable & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_consume;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_dout = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level != 5'd16);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_readable = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level != 1'd0);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_din = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_payload_data};
assign {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_payload_data} = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_ack = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_in_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_stb = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_eop = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_payload_data = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_fifo_out_payload_data;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_re = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_8;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr <= 4'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_replace) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_8 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_we = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_we & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_replace));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_do_read = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_readable & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_consume;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_dout = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level != 5'd16);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_readable = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level != 1'd0);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_trigger = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value != 1'd0);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_status;

// synthesis translate_off
reg dummy_d_9;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_clear <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_r)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_9 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_pending;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_irq = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_w & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_status = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_trigger;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_locked);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe = ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en[1] | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en[2]) | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en[3]);

// synthesis translate_off
reg dummy_d_10;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_valid <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_address <= 15'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_bank <= 3'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cke <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_odt <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_reset_n <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_mask <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_address <= 15'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_bank <= 3'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cke <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_odt <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_reset_n <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_mask <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_address <= 15'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_bank <= 3'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cke <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_odt <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_reset_n <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_mask <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_address <= 15'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_bank <= 3'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cke <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_odt <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_reset_n <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_mask <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_en <= 1'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[0]) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p0_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p1_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p2_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_slave_p3_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_valid;
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p0_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p1_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p2_rddata_valid;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_address;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_bank <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_bank;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cas_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cas_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_ras_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_ras_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_we_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_we_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_cke <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cke;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_odt <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_odt;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_reset_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_reset_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_wrdata_mask <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_mask;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_en <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_en;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_master_p3_rddata_valid;
	end
// synthesis translate_off
	dummy_d_10 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[1];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[1];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[1];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cke = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[1];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_odt = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[3];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[3];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[3];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_reset_n = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage[3];

// synthesis translate_off
reg dummy_d_11;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_we_n <= 1'd1;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cs_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[0]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_we_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[1]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cas_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[2]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_ras_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[3]);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cs_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_we_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_cas_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_11 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[4]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage[5]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_12;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_we_n <= 1'd1;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cs_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[0]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_we_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[1]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cas_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[2]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_ras_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[3]);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cs_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_we_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_cas_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_12 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[4]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage[5]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_13;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_we_n <= 1'd1;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cs_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[0]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_we_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[1]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cas_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[2]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_ras_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[3]);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cs_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_we_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_cas_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_13 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[4]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage[5]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_14;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_we_n <= 1'd1;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cs_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[0]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_we_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[1]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cas_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[2]);
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_ras_n <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[3]);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cs_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_we_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_cas_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_14 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_address = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[4]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_en = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_re & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage[5]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_wrdata_mask = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset1 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset2 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset3 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset4 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset5 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset6 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_open = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset7 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];

// synthesis translate_off
reg dummy_d_15;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7 <= 1'd0;
	case (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[9:7])
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0 <= 1'd1;
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1 <= 1'd1;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2 <= 1'd1;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3 <= 1'd1;
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4 <= 1'd1;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5 <= 1'd1;
		end
		3'd6: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6 <= 1'd1;
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_15 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_hit = ((((((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_hit & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_idle = ((((((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6)) | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_wait = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_wait = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_reset_n = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_odt = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cke = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cs_n = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_16;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address <= 15'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address <= 11'd1024;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
		end else begin
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read)) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_address <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_16 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_reset_n = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_odt = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cke = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cs_n = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_17;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address <= 15'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address <= 11'd1024;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
		end else begin
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read)) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_address <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_17 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_reset_n = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_odt = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cke = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cs_n = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_18;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address <= 15'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address <= 11'd1024;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
		end else begin
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read)) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_address <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_18 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_reset_n = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_odt = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cke = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_cs_n = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_bank = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_19;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address <= 15'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address <= 11'd1024;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[24:10];
		end else begin
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read)) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_address <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_19 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_r = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_rddata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_rddata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_rddata};
assign {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata} = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_w;
assign {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p3_wrdata_mask, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_mask, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_wrdata_mask, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_wrdata_mask} = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_sel);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_hit = ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row0 == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_done = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count == 1'd0);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_done = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count == 1'd0);

// synthesis translate_off
reg dummy_d_20;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cas_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_ras_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_we_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read <= 1'd0;
	minicon_next_state <= 6'd0;
	minicon_next_state <= minicon_state;
	case (minicon_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_read <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_en <= 1'd1;
			minicon_next_state <= 2'd2;
		end
		2'd2: begin
			if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_rddata_valid) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack <= 1'd1;
				minicon_next_state <= 1'd0;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_ras_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_cas_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_we_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p2_wrdata_en <= 1'd1;
			minicon_next_state <= 4'd9;
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack <= 1'd1;
			minicon_next_state <= 1'd0;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_precharge_all <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n <= 1'd0;
			minicon_next_state <= 4'd14;
		end
		3'd6: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_ras_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cas_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_we_n <= 1'd0;
			minicon_next_state <= 4'd10;
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_activate <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_ras_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_cas_n <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p0_we_n <= 1'd1;
			minicon_next_state <= 4'd12;
		end
		4'd8: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_ras_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_cas_n <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_dfi_p1_we_n <= 1'd1;
			minicon_next_state <= 5'd16;
		end
		4'd9: begin
			minicon_next_state <= 3'd4;
		end
		4'd10: begin
			minicon_next_state <= 4'd11;
		end
		4'd11: begin
			minicon_next_state <= 3'd7;
		end
		4'd12: begin
			minicon_next_state <= 4'd13;
		end
		4'd13: begin
			minicon_next_state <= 1'd0;
		end
		4'd14: begin
			minicon_next_state <= 4'd15;
		end
		4'd15: begin
			minicon_next_state <= 4'd8;
		end
		5'd16: begin
			minicon_next_state <= 5'd17;
		end
		5'd17: begin
			minicon_next_state <= 5'd18;
		end
		5'd18: begin
			minicon_next_state <= 5'd19;
		end
		5'd19: begin
			minicon_next_state <= 5'd20;
		end
		5'd20: begin
			minicon_next_state <= 5'd21;
		end
		5'd21: begin
			minicon_next_state <= 5'd22;
		end
		5'd22: begin
			minicon_next_state <= 5'd23;
		end
		5'd23: begin
			minicon_next_state <= 5'd24;
		end
		5'd24: begin
			minicon_next_state <= 5'd25;
		end
		5'd25: begin
			minicon_next_state <= 5'd26;
		end
		5'd26: begin
			minicon_next_state <= 5'd27;
		end
		5'd27: begin
			minicon_next_state <= 5'd28;
		end
		5'd28: begin
			minicon_next_state <= 5'd29;
		end
		5'd29: begin
			minicon_next_state <= 5'd30;
		end
		5'd30: begin
			minicon_next_state <= 5'd31;
		end
		5'd31: begin
			minicon_next_state <= 6'd32;
		end
		6'd32: begin
			minicon_next_state <= 6'd33;
		end
		6'd33: begin
			minicon_next_state <= 6'd34;
		end
		6'd34: begin
			minicon_next_state <= 6'd35;
		end
		6'd35: begin
			minicon_next_state <= 6'd36;
		end
		6'd36: begin
			minicon_next_state <= 6'd37;
		end
		6'd37: begin
			minicon_next_state <= 6'd38;
		end
		6'd38: begin
			minicon_next_state <= 6'd39;
		end
		6'd39: begin
			minicon_next_state <= 6'd40;
		end
		6'd40: begin
			minicon_next_state <= 6'd41;
		end
		6'd41: begin
			minicon_next_state <= 6'd42;
		end
		6'd42: begin
			minicon_next_state <= 6'd43;
		end
		6'd43: begin
			minicon_next_state <= 6'd44;
		end
		6'd44: begin
			minicon_next_state <= 6'd45;
		end
		6'd45: begin
			minicon_next_state <= 1'd0;
		end
		default: begin
			if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_done) begin
				minicon_next_state <= 3'd5;
			end else begin
				if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_stb & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_cyc)) begin
					if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_hit) begin
						if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_we) begin
							minicon_next_state <= 2'd3;
						end else begin
							minicon_next_state <= 1'd1;
						end
					end else begin
						if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank_idle)) begin
							if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_done) begin
								minicon_next_state <= 3'd6;
							end
						end else begin
							minicon_next_state <= 3'd7;
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_20 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[14:2];

// synthesis translate_off
reg dummy_d_21;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we <= 16'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w <= 128'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_write_from_slave) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_r;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we <= {16{1'd1}};
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w <= {4{monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_w}};
		if ((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_stb) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_we) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we <= {({4{(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[1:0] == 1'd0)}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel), ({4{(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[1:0] == 1'd1)}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel), ({4{(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[1:0] == 2'd2)}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel), ({4{(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[1:0] == 2'd3)}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel)};
		end
	end
// synthesis translate_off
	dummy_d_21 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_sel = 16'd65535;

// synthesis translate_off
reg dummy_d_22;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r <= 32'd0;
	case (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_adr_offset_r)
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[127:96];
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[95:64];
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[63:32];
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[31:0];
		end
	endcase
// synthesis translate_off
	dummy_d_22 <= dummy_s;
// synthesis translate_on
end
assign {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_dirty, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_tag} = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_w = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_dirty, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_tag};
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[14:2];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_tag = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[29:15];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_adr = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_tag, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[14:2]};

// synthesis translate_off
reg dummy_d_23;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_write_from_slave <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_dirty <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_clr <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_inc <= 1'd0;
	fullmemorywe_next_state <= 3'd0;
	fullmemorywe_next_state <= fullmemorywe_state;
	case (fullmemorywe_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_clr <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_tag == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[29:15])) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack <= 1'd1;
				if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_we) begin
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_di_dirty <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_we <= 1'd1;
				end
				fullmemorywe_next_state <= 1'd0;
			end else begin
				if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_do_dirty) begin
					fullmemorywe_next_state <= 2'd2;
				end else begin
					fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_we <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_ack) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_inc <= 1'd1;
				if (1'd1) begin
					fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_we <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_clr <= 1'd1;
			fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_we <= 1'd0;
			if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_ack) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_write_from_slave <= 1'd1;
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_word_inc <= 1'd1;
				if (1'd1) begin
					fullmemorywe_next_state <= 1'd1;
				end else begin
					fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_stb)) begin
				fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_23 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr;

// synthesis translate_off
reg dummy_d_24;
// synthesis translate_on
always @(*) begin
	spiflash2x_cs_n <= 1'd1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_status <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_o <= 2'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe <= 1'd0;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage[1];
		spiflash2x_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage[2];
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage[3]) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe <= 1'd0;
		end else begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe <= 1'd1;
		end
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage[1]) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i0[1];
		end
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_o <= {{1{1'd1}}, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage[0]};
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_clk;
		spiflash2x_cs_n <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_cs_n;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_o <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr[31:30];
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dq_oe;
	end
// synthesis translate_off
	dummy_d_24 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_reset = monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset0;
assign monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock0 = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_lock;
assign monroe_ionphoton_monroe_ionphoton_tx_reset = monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset0;
assign monroe_ionphoton_monroe_ionphoton_rx_init_enable = monroe_ionphoton_monroe_ionphoton_tx_init_done;
assign monroe_ionphoton_monroe_ionphoton_rx_reset = monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset0;
assign monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done0 = monroe_ionphoton_monroe_ionphoton_rx_pma_reset_done;
assign monroe_ionphoton_monroe_ionphoton_drpaddr = monroe_ionphoton_monroe_ionphoton_rx_init_drpaddr;
assign monroe_ionphoton_monroe_ionphoton_drpen = monroe_ionphoton_monroe_ionphoton_rx_init_drpen;
assign monroe_ionphoton_monroe_ionphoton_drpdi = monroe_ionphoton_monroe_ionphoton_rx_init_drpdi;
assign monroe_ionphoton_monroe_ionphoton_rx_init_drprdy = monroe_ionphoton_monroe_ionphoton_drprdy;
assign monroe_ionphoton_monroe_ionphoton_rx_init_drpdo = monroe_ionphoton_monroe_ionphoton_drpdo;
assign monroe_ionphoton_monroe_ionphoton_drpwe = monroe_ionphoton_monroe_ionphoton_rx_init_drpwe;
assign monroe_ionphoton_monroe_ionphoton_i = monroe_ionphoton_monroe_ionphoton_pcs_restart;
assign monroe_ionphoton_monroe_ionphoton_rx_init_restart = monroe_ionphoton_monroe_ionphoton_o;
assign monroe_ionphoton_monroe_ionphoton_tx_data0 = monroe_ionphoton_monroe_ionphoton_tx_data_half;
assign monroe_ionphoton_monroe_ionphoton_rx_data_half = monroe_ionphoton_monroe_ionphoton_rx_data0;
assign monroe_ionphoton_monroe_ionphoton_tx_data1 = monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output0;
assign monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input = monroe_ionphoton_monroe_ionphoton_rx_data1;
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_stb = monroe_ionphoton_monroe_ionphoton_pcs_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_ack = monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_ack;
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_data = monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_pcs_source_eop = ((~monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en) & monroe_ionphoton_monroe_ionphoton_pcs_rx_en_d);
assign monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_i = monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_valid_ci;
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg = (6'd32 | (monroe_ionphoton_monroe_ionphoton_pcs_autoneg_ack <<< 4'd14));
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1 = monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0;
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k1 = monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0;
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter = (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_in ^ monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_unbalanced);

// synthesis translate_off
reg dummy_d_25;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_6b <= 6'd0;
	if (((~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_in) & monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_flip)) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_6b <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b);
	end else begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_6b <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b;
	end
// synthesis translate_off
	dummy_d_25 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_26;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b <= 4'd0;
	if (((~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter) & monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0)) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter);
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b <= 3'd7;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter & monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1)) begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter);
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b <= 4'd8;
		end else begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out <= (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter ^ monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_unbalanced);
			if (((~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_inter) & monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_flip)) begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b);
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b;
			end
		end
	end
// synthesis translate_off
	dummy_d_26 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first = {monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_6b, monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_4b};

// synthesis translate_off
reg dummy_d_27;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1 <= 10'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[0] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[9];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[1] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[8];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[2] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[7];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[3] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[6];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[4] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[5];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[5] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[4];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[6] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[3];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[7] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[2];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[8] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[1];
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1[9] <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output_msb_first[0];
// synthesis translate_off
	dummy_d_27 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_28;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_load_config_reg_buffer <= 1'd0;
	a7_1000basex_transmitpath_next_state <= 3'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd0;
	a7_1000basex_transmitpath_next_state <= a7_1000basex_transmitpath_state;
	case (a7_1000basex_transmitpath_state)
		1'd1: begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type) begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 7'd66;
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd181;
			end
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type);
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value_ce <= 1'd1;
			a7_1000basex_transmitpath_next_state <= 2'd2;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg_buffer[7:0];
			a7_1000basex_transmitpath_next_state <= 2'd3;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg_buffer[15:8];
			a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd4: begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disparity) begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd197;
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 7'd80;
			end
			a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_ack <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_stb) begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_data;
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd253;
				a7_1000basex_transmitpath_next_state <= 3'd6;
			end
		end
		3'd6: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd247;
			if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_parity) begin
				a7_1000basex_transmitpath_next_state <= 1'd0;
			end else begin
				a7_1000basex_transmitpath_next_state <= 3'd7;
			end
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd247;
			a7_1000basex_transmitpath_next_state <= 1'd0;
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_ack <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb) begin
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_load_config_reg_buffer <= 1'd1;
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
				monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd188;
				a7_1000basex_transmitpath_next_state <= 1'd1;
			end else begin
				if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_tx_stb) begin
					monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd251;
					a7_1000basex_transmitpath_next_state <= 3'd5;
				end else begin
					monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k0 <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d0 <= 8'd188;
					a7_1000basex_transmitpath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_28 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_data = (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_first_preamble_byte ? 7'd85 : monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d);

// synthesis translate_off
reg dummy_d_29;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first <= 10'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[0] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[9];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[1] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[8];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[2] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[7];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[6];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[4] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[5];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[5] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[4];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[6] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[3];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[7] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[2];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[8] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[1];
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9] <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input[0];
// synthesis translate_off
	dummy_d_29 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d = {monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b, monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code5b};

// synthesis translate_off
reg dummy_d_30;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_valid_ci <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_lsb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_msb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_first_preamble_byte <= 1'd0;
	a7_1000basex_receivepath_next_state <= 3'd0;
	a7_1000basex_receivepath_next_state <= a7_1000basex_receivepath_state;
	case (a7_1000basex_receivepath_state)
		1'd1: begin
			a7_1000basex_receivepath_next_state <= 1'd0;
			if ((~monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k)) begin
				if (((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 8'd181) | (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 7'd66))) begin
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_valid_ci <= 1'd1;
					a7_1000basex_receivepath_next_state <= 2'd2;
				end
				if (((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 8'd197) | (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 7'd80))) begin
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_valid_ci <= 1'd1;
					a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end
		end
		2'd2: begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k) begin
				if ((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 8'd251)) begin
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_first_preamble_byte <= 1'd1;
					a7_1000basex_receivepath_next_state <= 3'd4;
				end else begin
					a7_1000basex_receivepath_next_state <= 1'd0;
				end
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_lsb <= 1'd1;
				a7_1000basex_receivepath_next_state <= 2'd3;
			end
		end
		2'd3: begin
			if ((~monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k)) begin
				monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_msb <= 1'd1;
			end
			a7_1000basex_receivepath_next_state <= 1'd0;
		end
		3'd4: begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k) begin
				a7_1000basex_receivepath_next_state <= 1'd0;
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en <= 1'd1;
			end
		end
		default: begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k) begin
				if ((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 8'd188)) begin
					a7_1000basex_receivepath_next_state <= 1'd1;
				end
				if ((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d == 8'd251)) begin
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_first_preamble_byte <= 1'd1;
					a7_1000basex_receivepath_next_state <= 3'd4;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_30 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_o = (monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o ^ monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_o = (monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o ^ monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_o = (monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o ^ monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_pcs_done = (monroe_ionphoton_monroe_ionphoton_pcs_count == 1'd0);

// synthesis translate_off
reg dummy_d_31;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_link_up <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_restart <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_autoneg_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_wait <= 1'd0;
	a7_1000basex_fsm_next_state <= 2'd0;
	a7_1000basex_fsm_next_state <= a7_1000basex_fsm_state;
	case (a7_1000basex_fsm_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_autoneg_ack <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_o) begin
				a7_1000basex_fsm_next_state <= 2'd2;
			end
			if ((monroe_ionphoton_monroe_ionphoton_pcs_checker_tick & (~monroe_ionphoton_monroe_ionphoton_pcs_checker_ok))) begin
				monroe_ionphoton_monroe_ionphoton_pcs_restart <= 1'd1;
				a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_autoneg_ack <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_wait <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_pcs_done) begin
				a7_1000basex_fsm_next_state <= 2'd3;
			end
			if ((monroe_ionphoton_monroe_ionphoton_pcs_checker_tick & (~monroe_ionphoton_monroe_ionphoton_pcs_checker_ok))) begin
				monroe_ionphoton_monroe_ionphoton_pcs_restart <= 1'd1;
				a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_pcs_link_up <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_pcs_checker_tick & (~monroe_ionphoton_monroe_ionphoton_pcs_checker_ok))) begin
				monroe_ionphoton_monroe_ionphoton_pcs_restart <= 1'd1;
				a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_stb <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_o | monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_o)) begin
				a7_1000basex_fsm_next_state <= 1'd1;
			end
			if ((monroe_ionphoton_monroe_ionphoton_pcs_checker_tick & (~monroe_ionphoton_monroe_ionphoton_pcs_checker_ok))) begin
				monroe_ionphoton_monroe_ionphoton_pcs_restart <= 1'd1;
				a7_1000basex_fsm_next_state <= 1'd0;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_31 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_32;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_init_done <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset1 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset1 <= 1'd0;
	a7_1000basex_gtptxinit_next_state <= 2'd0;
	a7_1000basex_gtptxinit_next_state <= a7_1000basex_gtptxinit_state;
	case (a7_1000basex_gtptxinit_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset1 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset1 <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_tx_init_tick) begin
				a7_1000basex_gtptxinit_next_state <= 2'd2;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset1 <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock1 & monroe_ionphoton_monroe_ionphoton_tx_init_tick)) begin
				a7_1000basex_gtptxinit_next_state <= 2'd3;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_tx_init_done <= 1'd1;
		end
		default: begin
			if (monroe_ionphoton_monroe_ionphoton_tx_init_tick) begin
				a7_1000basex_gtptxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_32 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_rx_init_drpaddr = 5'd17;

// synthesis translate_off
reg dummy_d_33;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_init_drpdi <= 16'd0;
	if (monroe_ionphoton_monroe_ionphoton_rx_init_drpmask) begin
		monroe_ionphoton_monroe_ionphoton_rx_init_drpdi <= (monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue & 16'd63487);
	end else begin
		monroe_ionphoton_monroe_ionphoton_rx_init_drpdi <= monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue;
	end
// synthesis translate_off
	dummy_d_33 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_34;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_init_drpen <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_drpwe <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_done <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_drpmask <= 1'd0;
	a7_1000basex_gtprxinit_next_state <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value <= 16'd0;
	monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd0;
	a7_1000basex_gtprxinit_next_state <= a7_1000basex_gtprxinit_state;
	case (a7_1000basex_gtprxinit_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd1;
			a7_1000basex_gtprxinit_next_state <= 2'd2;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_rx_init_drpen <= 1'd1;
			a7_1000basex_gtprxinit_next_state <= 2'd3;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_rx_init_drprdy) begin
				monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value <= monroe_ionphoton_monroe_ionphoton_rx_init_drpdo;
				monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value_ce <= 1'd1;
				a7_1000basex_gtprxinit_next_state <= 3'd4;
			end
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_rx_init_drpmask <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_rx_init_drpen <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_rx_init_drpwe <= 1'd1;
			a7_1000basex_gtprxinit_next_state <= 3'd5;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1 <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_rx_init_drprdy) begin
				a7_1000basex_gtprxinit_next_state <= 3'd6;
			end
		end
		3'd6: begin
			if ((monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done_r & (~monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done1))) begin
				a7_1000basex_gtprxinit_next_state <= 3'd7;
			end
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_drpen <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_rx_init_drpwe <= 1'd1;
			a7_1000basex_gtprxinit_next_state <= 4'd8;
		end
		4'd8: begin
			if (monroe_ionphoton_monroe_ionphoton_rx_init_drprdy) begin
				a7_1000basex_gtprxinit_next_state <= 4'd9;
			end
		end
		4'd9: begin
			monroe_ionphoton_monroe_ionphoton_rx_init_done <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_rx_init_restart) begin
				a7_1000basex_gtprxinit_next_state <= 1'd0;
			end
		end
		default: begin
			if (monroe_ionphoton_monroe_ionphoton_rx_init_enable) begin
				a7_1000basex_gtprxinit_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_34 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_o = (monroe_ionphoton_monroe_ionphoton_toggle_o ^ monroe_ionphoton_monroe_ionphoton_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_stb = monroe_ionphoton_monroe_ionphoton_source_stb;
assign monroe_ionphoton_monroe_ionphoton_source_ack = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_eop = monroe_ionphoton_monroe_ionphoton_source_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_data = monroe_ionphoton_monroe_ionphoton_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_error = monroe_ionphoton_monroe_ionphoton_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_sink_stb = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_ack = monroe_ionphoton_monroe_ionphoton_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_sink_eop = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_eop;
assign monroe_ionphoton_monroe_ionphoton_sink_payload_data = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_sink_payload_error = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_ps_preamble_error_i = monroe_ionphoton_monroe_ionphoton_preamble_checker_error;
assign monroe_ionphoton_monroe_ionphoton_ps_crc_error_i = monroe_ionphoton_monroe_ionphoton_crc32_checker_error;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_stb = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_ack = monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_eop = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_stb = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_ack = monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_eop = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_data = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_error = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_stb = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_source_ack = monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_eop = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_eop;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_data = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_error = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb = monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_source_ack = monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_eop = monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_data = monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_error = monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_stb = monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack = monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_eop = monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_error = monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_stb = monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_eop = monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_data = monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_error = monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_stb = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_ack = monroe_ionphoton_monroe_ionphoton_pcs_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_eop = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_data = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_pcs_sink_payload_error = monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_stb = monroe_ionphoton_monroe_ionphoton_pcs_source_stb;
assign monroe_ionphoton_monroe_ionphoton_pcs_source_ack = monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_eop = monroe_ionphoton_monroe_ionphoton_pcs_source_eop;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_data = monroe_ionphoton_monroe_ionphoton_pcs_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_pcs_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_error = monroe_ionphoton_monroe_ionphoton_pcs_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb = monroe_ionphoton_monroe_ionphoton_preamble_checker_source_stb;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_source_ack = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_eop = monroe_ionphoton_monroe_ionphoton_preamble_checker_source_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_data = monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_error = monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_stb = monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_stb;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_ack = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_eop = monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_eop;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_error = monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_stb = monroe_ionphoton_monroe_ionphoton_padding_checker_source_stb;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_ack = monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_eop = monroe_ionphoton_monroe_ionphoton_padding_checker_source_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_data = monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_error = monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_stb = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_source_ack = monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_eop = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_data = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_error = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_error;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_stb = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_ack = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_eop = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_data = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_error = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error;

// synthesis translate_off
reg dummy_d_35;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_data <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_last_be <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_ce <= 1'd0;
	liteethmacgap_next_state <= 1'd0;
	liteethmacgap_next_state <= liteethmacgap_state;
	case (liteethmacgap_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_ce <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter == 4'd11)) begin
				liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_reset <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_stb <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_stb;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_ack <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_ack;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_eop <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_eop;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_data;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_last_be <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_last_be;
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_source_payload_error <= monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_payload_error;
			if (((monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_stb & monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_eop) & monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_sink_ack)) begin
				liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_35 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_36;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_clr_cnt <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_inc_cnt <= 1'd0;
	liteethmacpreambleinserter_next_state <= 2'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_data;
	liteethmacpreambleinserter_next_state <= liteethmacpreambleinserter_state;
	case (liteethmacpreambleinserter_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_stb <= 1'd1;
			case (monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt)
				1'd0: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[55:48];
				end
				default: begin
					monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt == 3'd7)) begin
				if (monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack) begin
					liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				monroe_ionphoton_monroe_ionphoton_preamble_inserter_inc_cnt <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_stb <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_stb;
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack;
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_eop <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_eop;
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_payload_error <= monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_payload_error;
			if (((monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_stb & monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_eop) & monroe_ionphoton_monroe_ionphoton_preamble_inserter_source_ack)) begin
				liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_clr_cnt <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_stb) begin
				monroe_ionphoton_monroe_ionphoton_preamble_inserter_sink_ack <= 1'd0;
				liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_36 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_data = monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_37;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_checker_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_checker_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_preamble_checker_error <= 1'd0;
	liteethmacpreamblechecker_next_state <= 1'd0;
	liteethmacpreamblechecker_next_state <= liteethmacpreamblechecker_state;
	case (liteethmacpreamblechecker_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_preamble_checker_source_stb <= monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_stb;
			monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_ack <= monroe_ionphoton_monroe_ionphoton_preamble_checker_source_ack;
			monroe_ionphoton_monroe_ionphoton_preamble_checker_source_eop <= monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_eop;
			monroe_ionphoton_monroe_ionphoton_preamble_checker_source_payload_error <= monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_error;
			if (((monroe_ionphoton_monroe_ionphoton_preamble_checker_source_stb & monroe_ionphoton_monroe_ionphoton_preamble_checker_source_eop) & monroe_ionphoton_monroe_ionphoton_preamble_checker_source_ack)) begin
				liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_ack <= 1'd1;
			if (((monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_stb & (~monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_eop)) & (monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_payload_data == 8'd213))) begin
				liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_stb & monroe_ionphoton_monroe_ionphoton_preamble_checker_sink_eop)) begin
				monroe_ionphoton_monroe_ionphoton_preamble_checker_error <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_37 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt_done = (monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt == 1'd0);
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1 = monroe_ionphoton_monroe_ionphoton_crc32_inserter_data0;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_last = monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg;
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_value = (~{monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[0], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[1], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[2], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[3], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[4], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[5], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[6], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[7], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[8], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[9], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[10], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[11], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[12], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[13], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[14], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[15], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[16], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[17], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[18], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[19], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[20], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[21], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[22], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[23], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[24], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[25], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[26], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[27], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[28], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[29], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[30], monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg[31]});
assign monroe_ionphoton_monroe_ionphoton_crc32_inserter_error = (monroe_ionphoton_monroe_ionphoton_crc32_inserter_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_38;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[0] <= (((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[1] <= (((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[2] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[3] <= (((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[4] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[5] <= (((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[6] <= (((((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[7] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[8] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[0] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[9] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[1] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[10] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[2] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[11] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[3] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[12] <= ((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[4] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[13] <= ((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[5] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[14] <= ((((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[6] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[15] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[7] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[16] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[8] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[17] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[9] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[18] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[10] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[19] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[11] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[20] <= ((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[12] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[21] <= ((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[13] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[22] <= ((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[14] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[23] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[15] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[24] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[16] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[25] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[17] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[26] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[18] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[27] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[19] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[28] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[20] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[29] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[21] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[30] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[22] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[3]);
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_next[31] <= ((monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[23] ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_inserter_data1[2]);
// synthesis translate_off
	dummy_d_38 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_39;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_last_be <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_data0 <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_ce <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing0 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing1 <= 1'd0;
	liteethmaccrc32inserter_next_state <= 2'd0;
	liteethmaccrc32inserter_next_state <= liteethmaccrc32inserter_state;
	case (liteethmaccrc32inserter_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_ce <= (monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb & monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack);
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_data0 <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_data;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_stb <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_eop;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_data;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_last_be <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_last_be;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_error <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_payload_error;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop <= 1'd0;
			if (((monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb & monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_eop) & monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack)) begin
				liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_stb <= 1'd1;
			case (monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt)
				1'd0: begin
					monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_value[31:24];
				end
				1'd1: begin
					monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_value[23:16];
				end
				2'd2: begin
					monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_value[15:8];
				end
				default: begin
					monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_value[7:0];
				end
			endcase
			if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt_done) begin
				monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_eop <= 1'd1;
				if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack) begin
					liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_reset <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_stb) begin
				monroe_ionphoton_monroe_ionphoton_crc32_inserter_sink_ack <= 1'd0;
				liteethmaccrc32inserter_next_state <= 1'd1;
			end
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_39 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_full = (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level == 3'd4);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_in = (monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb & ((~monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_full) | monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_out));
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_out = (monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_stb & monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_ack);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_eop = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_error = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_error;

// synthesis translate_off
reg dummy_d_40;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_stb <= monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_stb <= monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_40 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_41;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack <= monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_ack;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack <= monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_41 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_stb = (monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_full);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_eop = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_ack = monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_out;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_last_be;

// synthesis translate_off
reg dummy_d_42;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_error <= monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_error;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_payload_error <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_error | monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_error);
// synthesis translate_off
	dummy_d_42 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_error = ((monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_stb & monroe_ionphoton_monroe_ionphoton_crc32_checker_source_source_eop) & monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_error);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data0 = monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1 = monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data0;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last = monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_value = (~{monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[0], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[1], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[2], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[3], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[4], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[5], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[6], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[7], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[8], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[9], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[10], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[11], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[12], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[13], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[14], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[15], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[16], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[17], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[18], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[19], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[20], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[21], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[22], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[23], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[24], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[25], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[26], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[27], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[28], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[29], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[30], monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg[31]});
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_error = (monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_43;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[0] <= (((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[1] <= (((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[2] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[3] <= (((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[4] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[5] <= (((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[6] <= (((((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[7] <= (((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[8] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[0] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[9] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[1] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[10] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[2] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[11] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[3] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[12] <= ((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[4] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[13] <= ((((((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[5] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[14] <= ((((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[6] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[15] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[7] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[16] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[8] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[17] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[9] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[18] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[10] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[19] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[11] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[20] <= ((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[12] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[21] <= ((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[13] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[22] <= ((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[14] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[23] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[15] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[24] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[16] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[25] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[17] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[26] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[18] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[24]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[7]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[27] <= ((((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[19] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[25]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[6]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[28] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[20] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[26]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[5]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[29] <= ((((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[21] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[30]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[1]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[27]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[4]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[30] <= ((((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[22] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[31]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[0]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[28]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[3]);
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next[31] <= ((monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[23] ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_last[29]) ^ monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_data1[2]);
// synthesis translate_off
	dummy_d_43 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_din = {monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_error, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_last_be, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_data};
assign {monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_error, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_last_be, monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_data} = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_ack = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_we = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_in_payload_error = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_sink_payload_error;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_stb = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_eop = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_data = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_data;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_payload_error = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_fifo_out_payload_error;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_re = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_source_ack;

// synthesis translate_off
reg dummy_d_44;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_replace) begin
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr <= monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce;
	end
// synthesis translate_off
	dummy_d_44 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_we = (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_we & (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable | monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_replace));
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_do_read = (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_readable & monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_adr = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_dout = monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_dat_r;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable = (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level != 3'd5);
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_readable = (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_45;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_ce <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_reset <= 1'd0;
	liteethmaccrc32checker_next_state <= 2'd0;
	liteethmaccrc32checker_next_state <= liteethmaccrc32checker_state;
	case (liteethmaccrc32checker_state)
		1'd1: begin
			if ((monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack)) begin
				monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_ce <= 1'd1;
				liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_ack)) begin
				monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_ce <= 1'd1;
				if (monroe_ionphoton_monroe_ionphoton_crc32_checker_sink_sink_eop) begin
					liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reset <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_reset <= 1'd1;
			liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_45 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_ps_preamble_error_o = (monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o ^ monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_ps_crc_error_o = (monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o ^ monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o_r);
assign monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_done = (monroe_ionphoton_monroe_ionphoton_padding_inserter_counter >= 6'd59);

// synthesis translate_off
reg dummy_d_46;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_data <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_last_be <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_error <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_ce <= 1'd0;
	liteethmacpaddinginserter_next_state <= 1'd0;
	liteethmacpaddinginserter_next_state <= liteethmacpaddinginserter_state;
	case (liteethmacpaddinginserter_state)
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop <= monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_done;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_data <= 1'd0;
			if ((monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb & monroe_ionphoton_monroe_ionphoton_padding_inserter_source_ack)) begin
				monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_ce <= 1'd1;
				if (monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_done) begin
					monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_reset <= 1'd1;
					liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb <= monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_stb;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_ack <= monroe_ionphoton_monroe_ionphoton_padding_inserter_source_ack;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop <= monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_eop;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_data;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_last_be <= monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_last_be;
			monroe_ionphoton_monroe_ionphoton_padding_inserter_source_payload_error <= monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_payload_error;
			if ((monroe_ionphoton_monroe_ionphoton_padding_inserter_source_stb & monroe_ionphoton_monroe_ionphoton_padding_inserter_source_ack)) begin
				monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_ce <= 1'd1;
				if (monroe_ionphoton_monroe_ionphoton_padding_inserter_sink_eop) begin
					if ((~monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_done)) begin
						monroe_ionphoton_monroe_ionphoton_padding_inserter_source_eop <= 1'd0;
						liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_46 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_stb = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_sink_ack = monroe_ionphoton_monroe_ionphoton_padding_checker_source_ack;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_eop = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_data = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_padding_checker_source_payload_error = monroe_ionphoton_monroe_ionphoton_padding_checker_sink_payload_error;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_source_stb = (monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_stb & monroe_ionphoton_monroe_ionphoton_tx_last_be_ongoing);
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_source_eop = monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_source_payload_data = monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_ack = monroe_ionphoton_monroe_ionphoton_tx_last_be_source_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_source_stb = monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_ack = monroe_ionphoton_monroe_ionphoton_rx_last_be_source_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_source_eop = monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_data = monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_error = monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_error;

// synthesis translate_off
reg dummy_d_47;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_last_be <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_last_be <= monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_payload_last_be;
	monroe_ionphoton_monroe_ionphoton_rx_last_be_source_payload_last_be <= monroe_ionphoton_monroe_ionphoton_rx_last_be_sink_eop;
// synthesis translate_off
	dummy_d_47 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_stb = monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_eop = monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_ack = monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_ack;

// synthesis translate_off
reg dummy_d_48;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data <= 40'd0;
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[7:0] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data[7:0];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[8] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be[0];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[9] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error[0];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[17:10] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data[15:8];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[18] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be[1];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[19] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error[1];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[27:20] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data[23:16];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[28] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be[2];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[29] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error[2];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[37:30] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_data[31:24];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[38] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_last_be[3];
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[39] <= monroe_ionphoton_monroe_ionphoton_tx_converter_sink_sink_payload_error[3];
// synthesis translate_off
	dummy_d_48 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_stb = monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_eop = monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_ack = monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_ack;
assign {monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_error, monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_last_be, monroe_ionphoton_monroe_ionphoton_tx_converter_source_source_payload_data} = monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_last = (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux == 2'd3);
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_stb = monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_eop = (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_eop & monroe_ionphoton_monroe_ionphoton_tx_converter_converter_last);
assign monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_ack = (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_last & monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_ack);

// synthesis translate_off
reg dummy_d_49;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data <= 10'd0;
	case (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux)
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[39:30];
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[19:10];
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_payload_data <= monroe_ionphoton_monroe_ionphoton_tx_converter_converter_sink_payload_data[9:0];
		end
	endcase
// synthesis translate_off
	dummy_d_49 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_stb = monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_eop = monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_ack = monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data = {monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_error, monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_last_be, monroe_ionphoton_monroe_ionphoton_rx_converter_sink_sink_payload_data};
assign monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_stb = monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_eop = monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_ack = monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_ack;

// synthesis translate_off
reg dummy_d_50;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data[7:0] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[7:0];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data[15:8] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[17:10];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data[23:16] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[27:20];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_data[31:24] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[37:30];
// synthesis translate_off
	dummy_d_50 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_51;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be[0] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[8];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be[1] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[18];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be[2] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[28];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_last_be[3] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[38];
// synthesis translate_off
	dummy_d_51 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_52;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error[0] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[9];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error[1] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[19];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error[2] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[29];
	monroe_ionphoton_monroe_ionphoton_rx_converter_source_source_payload_error[3] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[39];
// synthesis translate_off
	dummy_d_52 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_ack = ((~monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all) | monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_ack);
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_stb = monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all;
assign monroe_ionphoton_monroe_ionphoton_rx_converter_converter_load_part = (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_stb & monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_ack);
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_din = {monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_error, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_last_be, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_data};
assign {monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_error, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_last_be, monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_data} = monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_ack = monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_we = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_data = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_in_payload_error = monroe_ionphoton_monroe_ionphoton_tx_cdc_sink_payload_error;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_stb = monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_eop = monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_data = monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_data;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_source_payload_error = monroe_ionphoton_monroe_ionphoton_tx_cdc_fifo_out_payload_error;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_re = monroe_ionphoton_monroe_ionphoton_tx_cdc_source_ack;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_ce = (monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_writable & monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_we);
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_ce = (monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_readable & monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_writable = (((monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q[6] == monroe_ionphoton_monroe_ionphoton_tx_cdc_consume_wdomain[6]) | (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q[5] == monroe_ionphoton_monroe_ionphoton_tx_cdc_consume_wdomain[5])) | (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q[4:0] != monroe_ionphoton_monroe_ionphoton_tx_cdc_consume_wdomain[4:0]));
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_readable = (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q != monroe_ionphoton_monroe_ionphoton_tx_cdc_produce_rdomain);
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_adr = monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary[5:0];
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_we = monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_ce;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_adr = monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary[5:0];
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_asyncfifo_dout = monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_53;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_ce) begin
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary <= (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_53 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next = (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary ^ monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_54;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_ce) begin
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary <= (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_54 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next = (monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary ^ monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary[6:1]);
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_din = {monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_error, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_last_be, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_data};
assign {monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_error, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_last_be, monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_data} = monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_ack = monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_we = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_data = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_last_be = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_in_payload_error = monroe_ionphoton_monroe_ionphoton_rx_cdc_sink_payload_error;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_stb = monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_eop = monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_data = monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_data;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_source_payload_error = monroe_ionphoton_monroe_ionphoton_rx_cdc_fifo_out_payload_error;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_re = monroe_ionphoton_monroe_ionphoton_rx_cdc_source_ack;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_ce = (monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_writable & monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_we);
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_ce = (monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_readable & monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_writable = (((monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q[6] == monroe_ionphoton_monroe_ionphoton_rx_cdc_consume_wdomain[6]) | (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q[5] == monroe_ionphoton_monroe_ionphoton_rx_cdc_consume_wdomain[5])) | (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q[4:0] != monroe_ionphoton_monroe_ionphoton_rx_cdc_consume_wdomain[4:0]));
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_readable = (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q != monroe_ionphoton_monroe_ionphoton_rx_cdc_produce_rdomain);
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_adr = monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary[5:0];
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_we = monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_ce;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_adr = monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary[5:0];
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_asyncfifo_dout = monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_55;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_ce) begin
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary <= (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_55 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next = (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary ^ monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_56;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_ce) begin
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary <= (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_56 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next = (monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary ^ monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary[6:1]);
assign monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb = monroe_ionphoton_monroe_ionphoton_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_sink_ack = monroe_ionphoton_monroe_ionphoton_writer_sink_sink_ack;
assign monroe_ionphoton_monroe_ionphoton_writer_sink_sink_eop = monroe_ionphoton_monroe_ionphoton_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data = monroe_ionphoton_monroe_ionphoton_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be = monroe_ionphoton_monroe_ionphoton_sink_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_error = monroe_ionphoton_monroe_ionphoton_sink_payload_error;
assign monroe_ionphoton_monroe_ionphoton_source_stb = monroe_ionphoton_monroe_ionphoton_reader_source_source_stb;
assign monroe_ionphoton_monroe_ionphoton_reader_source_source_ack = monroe_ionphoton_monroe_ionphoton_source_ack;
assign monroe_ionphoton_monroe_ionphoton_source_eop = monroe_ionphoton_monroe_ionphoton_reader_source_source_eop;
assign monroe_ionphoton_monroe_ionphoton_source_payload_data = monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data;
assign monroe_ionphoton_monroe_ionphoton_source_payload_last_be = monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be;
assign monroe_ionphoton_monroe_ionphoton_source_payload_error = monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_error;

// synthesis translate_off
reg dummy_d_57;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_writer_increment <= 3'd0;
	if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be[3]) begin
		monroe_ionphoton_monroe_ionphoton_writer_increment <= 1'd1;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be[2]) begin
			monroe_ionphoton_monroe_ionphoton_writer_increment <= 2'd2;
		end else begin
			if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be[1]) begin
				monroe_ionphoton_monroe_ionphoton_writer_increment <= 2'd3;
			end else begin
				monroe_ionphoton_monroe_ionphoton_writer_increment <= 3'd4;
			end
		end
	end
// synthesis translate_off
	dummy_d_57 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_slot = monroe_ionphoton_monroe_ionphoton_writer_slot;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_length = monroe_ionphoton_monroe_ionphoton_writer_counter;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_source_ack = monroe_ionphoton_monroe_ionphoton_writer_available_clear;
assign monroe_ionphoton_monroe_ionphoton_writer_available_trigger = monroe_ionphoton_monroe_ionphoton_writer_fifo_source_stb;
assign monroe_ionphoton_monroe_ionphoton_writer_slot_status = monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_slot;
assign monroe_ionphoton_monroe_ionphoton_writer_length_status = monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_length;

// synthesis translate_off
reg dummy_d_58;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_writer_memory0_adr <= 9'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory0_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_w <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory1_adr <= 9'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory1_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_w <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory2_adr <= 9'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory2_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_w <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory3_adr <= 9'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory3_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_w <= 32'd0;
	case (monroe_ionphoton_monroe_ionphoton_writer_slot)
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_writer_memory0_adr <= monroe_ionphoton_monroe_ionphoton_writer_counter[31:2];
			monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_w <= monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data;
			if ((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_writer_ongoing)) begin
				monroe_ionphoton_monroe_ionphoton_writer_memory0_we <= 4'd15;
			end
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_writer_memory1_adr <= monroe_ionphoton_monroe_ionphoton_writer_counter[31:2];
			monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_w <= monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data;
			if ((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_writer_ongoing)) begin
				monroe_ionphoton_monroe_ionphoton_writer_memory1_we <= 4'd15;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_writer_memory2_adr <= monroe_ionphoton_monroe_ionphoton_writer_counter[31:2];
			monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_w <= monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data;
			if ((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_writer_ongoing)) begin
				monroe_ionphoton_monroe_ionphoton_writer_memory2_we <= 4'd15;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_writer_memory3_adr <= monroe_ionphoton_monroe_ionphoton_writer_counter[31:2];
			monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_w <= monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_data;
			if ((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_writer_ongoing)) begin
				monroe_ionphoton_monroe_ionphoton_writer_memory3_we <= 4'd15;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_58 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_writer_status_w = monroe_ionphoton_monroe_ionphoton_writer_available_status;

// synthesis translate_off
reg dummy_d_59;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_writer_available_clear <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_writer_pending_re & monroe_ionphoton_monroe_ionphoton_writer_pending_r)) begin
		monroe_ionphoton_monroe_ionphoton_writer_available_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_59 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_writer_pending_w = monroe_ionphoton_monroe_ionphoton_writer_available_pending;
assign monroe_ionphoton_monroe_ionphoton_writer_irq = (monroe_ionphoton_monroe_ionphoton_writer_pending_w & monroe_ionphoton_monroe_ionphoton_writer_storage);
assign monroe_ionphoton_monroe_ionphoton_writer_available_status = monroe_ionphoton_monroe_ionphoton_writer_available_trigger;
assign monroe_ionphoton_monroe_ionphoton_writer_available_pending = monroe_ionphoton_monroe_ionphoton_writer_available_trigger;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_din = {monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_length, monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_slot};
assign {monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_length, monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_slot} = monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_ack = monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_we = monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_slot = monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_slot;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_in_payload_length = monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_payload_length;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_source_stb = monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_source_eop = monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_slot = monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_slot;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_source_payload_length = monroe_ionphoton_monroe_ionphoton_writer_fifo_fifo_out_payload_length;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_re = monroe_ionphoton_monroe_ionphoton_writer_fifo_source_ack;

// synthesis translate_off
reg dummy_d_60;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr <= 2'd0;
	if (monroe_ionphoton_monroe_ionphoton_writer_fifo_replace) begin
		monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr <= (monroe_ionphoton_monroe_ionphoton_writer_fifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr <= monroe_ionphoton_monroe_ionphoton_writer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_60 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_we = (monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_we & (monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable | monroe_ionphoton_monroe_ionphoton_writer_fifo_replace));
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_do_read = (monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_readable & monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_adr = monroe_ionphoton_monroe_ionphoton_writer_fifo_consume;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_dout = monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_dat_r;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable = (monroe_ionphoton_monroe_ionphoton_writer_fifo_level != 3'd4);
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_readable = (monroe_ionphoton_monroe_ionphoton_writer_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_61;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_writer_counter_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_counter_ce <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_slot_ce <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_ongoing <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_stb <= 1'd0;
	liteethmacsramwriter_next_state <= 2'd0;
	monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value <= 32'd0;
	monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value_ce <= 1'd0;
	liteethmacsramwriter_next_state <= liteethmacsramwriter_state;
	case (liteethmacsramwriter_state)
		1'd1: begin
			if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb) begin
				if ((monroe_ionphoton_monroe_ionphoton_writer_counter == 11'd1530)) begin
					liteethmacsramwriter_next_state <= 2'd2;
				end else begin
					monroe_ionphoton_monroe_ionphoton_writer_counter_ce <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_writer_ongoing <= 1'd1;
				end
				if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_eop) begin
					if (((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_error & monroe_ionphoton_monroe_ionphoton_writer_sink_sink_payload_last_be) != 1'd0)) begin
						monroe_ionphoton_monroe_ionphoton_writer_counter_reset <= 1'd1;
						liteethmacsramwriter_next_state <= 1'd0;
					end else begin
						liteethmacsramwriter_next_state <= 2'd3;
					end
				end
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_writer_counter_reset <= 1'd1;
			if ((monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb & monroe_ionphoton_monroe_ionphoton_writer_sink_sink_eop)) begin
				monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value <= (monroe_ionphoton_monroe_ionphoton_writer_errors_status + 1'd1);
				monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value_ce <= 1'd1;
				liteethmacsramwriter_next_state <= 1'd0;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_writer_counter_reset <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_writer_slot_ce <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_stb <= 1'd1;
			liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (monroe_ionphoton_monroe_ionphoton_writer_sink_sink_stb) begin
				if (monroe_ionphoton_monroe_ionphoton_writer_fifo_sink_ack) begin
					monroe_ionphoton_monroe_ionphoton_writer_ongoing <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_writer_counter_ce <= 1'd1;
					liteethmacsramwriter_next_state <= 1'd1;
				end else begin
					liteethmacsramwriter_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_61 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_stb = monroe_ionphoton_monroe_ionphoton_reader_start_re;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_slot = monroe_ionphoton_monroe_ionphoton_reader_slot_storage;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_length = monroe_ionphoton_monroe_ionphoton_reader_length_storage;
assign monroe_ionphoton_monroe_ionphoton_reader_ready_status = monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_ack;

// synthesis translate_off
reg dummy_d_62;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be <= 4'd0;
	if (monroe_ionphoton_monroe_ionphoton_reader_last) begin
		if ((monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length[1:0] == 2'd3)) begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be <= 2'd2;
		end else begin
			if ((monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length[1:0] == 2'd2)) begin
				monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be <= 3'd4;
			end else begin
				if ((monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length[1:0] == 1'd1)) begin
					monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be <= 4'd8;
				end else begin
					monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_last_be <= 1'd1;
				end
			end
		end
	end
// synthesis translate_off
	dummy_d_62 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_reader_last = ((monroe_ionphoton_monroe_ionphoton_reader_counter + 3'd4) >= monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length);
assign monroe_ionphoton_monroe_ionphoton_reader_memory0_adr = monroe_ionphoton_monroe_ionphoton_reader_counter[10:2];
assign monroe_ionphoton_monroe_ionphoton_reader_memory1_adr = monroe_ionphoton_monroe_ionphoton_reader_counter[10:2];
assign monroe_ionphoton_monroe_ionphoton_reader_memory2_adr = monroe_ionphoton_monroe_ionphoton_reader_counter[10:2];
assign monroe_ionphoton_monroe_ionphoton_reader_memory3_adr = monroe_ionphoton_monroe_ionphoton_reader_counter[10:2];

// synthesis translate_off
reg dummy_d_63;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data <= 32'd0;
	case (monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_slot)
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data <= monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r;
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data <= monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data <= monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_payload_data <= monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r;
		end
	endcase
// synthesis translate_off
	dummy_d_63 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_w = monroe_ionphoton_monroe_ionphoton_reader_done_status;

// synthesis translate_off
reg dummy_d_64;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_reader_done_clear <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_re & monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_r)) begin
		monroe_ionphoton_monroe_ionphoton_reader_done_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_64 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_w = monroe_ionphoton_monroe_ionphoton_reader_done_pending;
assign monroe_ionphoton_monroe_ionphoton_reader_irq = (monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_w & monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage);
assign monroe_ionphoton_monroe_ionphoton_reader_done_status = 1'd0;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_din = {monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_eop, monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_length, monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_slot};
assign {monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_eop, monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_length, monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_slot} = monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_dout;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_ack = monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_we = monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_eop = monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_eop;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_slot = monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_slot;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_in_payload_length = monroe_ionphoton_monroe_ionphoton_reader_fifo_sink_payload_length;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_source_stb = monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_readable;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_source_eop = monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_eop;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_slot = monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_slot;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_source_payload_length = monroe_ionphoton_monroe_ionphoton_reader_fifo_fifo_out_payload_length;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_re = monroe_ionphoton_monroe_ionphoton_reader_fifo_source_ack;

// synthesis translate_off
reg dummy_d_65;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr <= 2'd0;
	if (monroe_ionphoton_monroe_ionphoton_reader_fifo_replace) begin
		monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr <= (monroe_ionphoton_monroe_ionphoton_reader_fifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr <= monroe_ionphoton_monroe_ionphoton_reader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_65 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_dat_w = monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_din;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_we = (monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_we & (monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable | monroe_ionphoton_monroe_ionphoton_reader_fifo_replace));
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_do_read = (monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_readable & monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_re);
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_adr = monroe_ionphoton_monroe_ionphoton_reader_fifo_consume;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_dout = monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_dat_r;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable = (monroe_ionphoton_monroe_ionphoton_reader_fifo_level != 3'd4);
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_readable = (monroe_ionphoton_monroe_ionphoton_reader_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_66;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_reader_source_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_reader_source_source_eop <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_reader_done_trigger <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_reader_fifo_source_ack <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_reader_counter_reset <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_reader_counter_ce <= 1'd0;
	liteethmacsramreader_next_state <= 2'd0;
	liteethmacsramreader_next_state <= liteethmacsramreader_state;
	case (liteethmacsramreader_state)
		1'd1: begin
			if ((~monroe_ionphoton_monroe_ionphoton_reader_last_d)) begin
				liteethmacsramreader_next_state <= 2'd2;
			end else begin
				liteethmacsramreader_next_state <= 2'd3;
			end
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_reader_source_source_stb <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_reader_source_source_eop <= monroe_ionphoton_monroe_ionphoton_reader_last;
			if (monroe_ionphoton_monroe_ionphoton_reader_source_source_ack) begin
				monroe_ionphoton_monroe_ionphoton_reader_counter_ce <= (~monroe_ionphoton_monroe_ionphoton_reader_last);
				liteethmacsramreader_next_state <= 1'd1;
			end
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_reader_fifo_source_ack <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_reader_done_trigger <= 1'd1;
			liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			monroe_ionphoton_monroe_ionphoton_reader_counter_reset <= 1'd1;
			if (monroe_ionphoton_monroe_ionphoton_reader_fifo_source_stb) begin
				liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_66 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_ev_irq = (monroe_ionphoton_monroe_ionphoton_writer_irq | monroe_ionphoton_monroe_ionphoton_reader_irq);
assign monroe_ionphoton_monroe_ionphoton_sram0_adr0 = monroe_ionphoton_monroe_ionphoton_sram0_bus_adr0[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r0 = monroe_ionphoton_monroe_ionphoton_sram0_dat_r0;
assign monroe_ionphoton_monroe_ionphoton_sram1_adr0 = monroe_ionphoton_monroe_ionphoton_sram1_bus_adr0[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r0 = monroe_ionphoton_monroe_ionphoton_sram1_dat_r0;
assign monroe_ionphoton_monroe_ionphoton_sram2_adr0 = monroe_ionphoton_monroe_ionphoton_sram2_bus_adr0[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r0 = monroe_ionphoton_monroe_ionphoton_sram2_dat_r0;
assign monroe_ionphoton_monroe_ionphoton_sram3_adr0 = monroe_ionphoton_monroe_ionphoton_sram3_bus_adr0[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r0 = monroe_ionphoton_monroe_ionphoton_sram3_dat_r0;

// synthesis translate_off
reg dummy_d_67;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_sram0_we <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_sram0_we[0] <= (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1[0]);
	monroe_ionphoton_monroe_ionphoton_sram0_we[1] <= (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1[1]);
	monroe_ionphoton_monroe_ionphoton_sram0_we[2] <= (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1[2]);
	monroe_ionphoton_monroe_ionphoton_sram0_we[3] <= (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1[3]);
// synthesis translate_off
	dummy_d_67 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_sram0_adr1 = monroe_ionphoton_monroe_ionphoton_sram0_bus_adr1[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r1 = monroe_ionphoton_monroe_ionphoton_sram0_dat_r1;
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_w = monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_w1;

// synthesis translate_off
reg dummy_d_68;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_sram1_we <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_sram1_we[0] <= (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1[0]);
	monroe_ionphoton_monroe_ionphoton_sram1_we[1] <= (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1[1]);
	monroe_ionphoton_monroe_ionphoton_sram1_we[2] <= (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1[2]);
	monroe_ionphoton_monroe_ionphoton_sram1_we[3] <= (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1[3]);
// synthesis translate_off
	dummy_d_68 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_sram1_adr1 = monroe_ionphoton_monroe_ionphoton_sram1_bus_adr1[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r1 = monroe_ionphoton_monroe_ionphoton_sram1_dat_r1;
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_w = monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_w1;

// synthesis translate_off
reg dummy_d_69;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_sram2_we <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_sram2_we[0] <= (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1[0]);
	monroe_ionphoton_monroe_ionphoton_sram2_we[1] <= (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1[1]);
	monroe_ionphoton_monroe_ionphoton_sram2_we[2] <= (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1[2]);
	monroe_ionphoton_monroe_ionphoton_sram2_we[3] <= (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1[3]);
// synthesis translate_off
	dummy_d_69 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_sram2_adr1 = monroe_ionphoton_monroe_ionphoton_sram2_bus_adr1[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r1 = monroe_ionphoton_monroe_ionphoton_sram2_dat_r1;
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_w = monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_w1;

// synthesis translate_off
reg dummy_d_70;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_sram3_we <= 4'd0;
	monroe_ionphoton_monroe_ionphoton_sram3_we[0] <= (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1[0]);
	monroe_ionphoton_monroe_ionphoton_sram3_we[1] <= (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1[1]);
	monroe_ionphoton_monroe_ionphoton_sram3_we[2] <= (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1[2]);
	monroe_ionphoton_monroe_ionphoton_sram3_we[3] <= (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_we1) & monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1[3]);
// synthesis translate_off
	dummy_d_70 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_sram3_adr1 = monroe_ionphoton_monroe_ionphoton_sram3_bus_adr1[8:0];
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r1 = monroe_ionphoton_monroe_ionphoton_sram3_dat_r1;
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_w = monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_w1;

// synthesis translate_off
reg dummy_d_71;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_monroe_ionphoton_slave_sel <= 8'd0;
	monroe_ionphoton_monroe_ionphoton_slave_sel[0] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 1'd0);
	monroe_ionphoton_monroe_ionphoton_slave_sel[1] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 1'd1);
	monroe_ionphoton_monroe_ionphoton_slave_sel[2] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 2'd2);
	monroe_ionphoton_monroe_ionphoton_slave_sel[3] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 2'd3);
	monroe_ionphoton_monroe_ionphoton_slave_sel[4] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 3'd4);
	monroe_ionphoton_monroe_ionphoton_slave_sel[5] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 3'd5);
	monroe_ionphoton_monroe_ionphoton_slave_sel[6] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 3'd6);
	monroe_ionphoton_monroe_ionphoton_slave_sel[7] <= (monroe_ionphoton_monroe_ionphoton_bus_adr[11:9] == 3'd7);
// synthesis translate_off
	dummy_d_71 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_adr0 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_w0 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_sel0 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_stb0 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_we0 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_cti0 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_bte0 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_adr0 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_w0 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_sel0 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_stb0 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_we0 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_cti0 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_bte0 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_adr0 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_w0 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_sel0 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_stb0 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_we0 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_cti0 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_bte0 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_adr0 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_w0 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_sel0 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_stb0 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_we0 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_cti0 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_bte0 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_adr1 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_w1 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_sel1 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_we1 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_cti1 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_bte1 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_adr1 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_w1 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_sel1 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_we1 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_cti1 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_bte1 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_adr1 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_w1 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_sel1 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_we1 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_cti1 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_bte1 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_adr1 = monroe_ionphoton_monroe_ionphoton_bus_adr;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_w1 = monroe_ionphoton_monroe_ionphoton_bus_dat_w;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_sel1 = monroe_ionphoton_monroe_ionphoton_bus_sel;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1 = monroe_ionphoton_monroe_ionphoton_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_we1 = monroe_ionphoton_monroe_ionphoton_bus_we;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_cti1 = monroe_ionphoton_monroe_ionphoton_bus_cti;
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_bte1 = monroe_ionphoton_monroe_ionphoton_bus_bte;
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc0 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[0]);
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc0 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[1]);
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc0 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[2]);
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc0 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[3]);
assign monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[4]);
assign monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[5]);
assign monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[6]);
assign monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 = (monroe_ionphoton_monroe_ionphoton_bus_cyc & monroe_ionphoton_monroe_ionphoton_slave_sel[7]);
assign monroe_ionphoton_monroe_ionphoton_bus_ack = (((((((monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0 | monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0) | monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0) | monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0) | monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1) | monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1) | monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1) | monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1);
assign monroe_ionphoton_monroe_ionphoton_bus_err = (((((((monroe_ionphoton_monroe_ionphoton_sram0_bus_err0 | monroe_ionphoton_monroe_ionphoton_sram1_bus_err0) | monroe_ionphoton_monroe_ionphoton_sram2_bus_err0) | monroe_ionphoton_monroe_ionphoton_sram3_bus_err0) | monroe_ionphoton_monroe_ionphoton_sram0_bus_err1) | monroe_ionphoton_monroe_ionphoton_sram1_bus_err1) | monroe_ionphoton_monroe_ionphoton_sram2_bus_err1) | monroe_ionphoton_monroe_ionphoton_sram3_bus_err1);
assign monroe_ionphoton_monroe_ionphoton_bus_dat_r = (((((((({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[0]}} & monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r0) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[1]}} & monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r0)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[2]}} & monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r0)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[3]}} & monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r0)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[4]}} & monroe_ionphoton_monroe_ionphoton_sram0_bus_dat_r1)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[5]}} & monroe_ionphoton_monroe_ionphoton_sram1_bus_dat_r1)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[6]}} & monroe_ionphoton_monroe_ionphoton_sram2_bus_dat_r1)) | ({32{monroe_ionphoton_monroe_ionphoton_slave_sel_r[7]}} & monroe_ionphoton_monroe_ionphoton_sram3_bus_dat_r1));
assign sys_kernel_clk = sys_clk;
assign sys_kernel_rst = monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_adr = monroe_ionphoton_monroe_ionphoton_kernel_cpu_i_adr_o[31:2];
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_adr = monroe_ionphoton_monroe_ionphoton_kernel_cpu_d_adr_o[31:2];
assign shared_adr = comb_rhs_array_muxed0;
assign shared_dat_w = comb_rhs_array_muxed1;
assign shared_sel = comb_rhs_array_muxed2;
assign shared_cyc = comb_rhs_array_muxed3;
assign shared_stb = comb_rhs_array_muxed4;
assign shared_we = comb_rhs_array_muxed5;
assign shared_cti = comb_rhs_array_muxed6;
assign shared_bte = comb_rhs_array_muxed7;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_r = shared_dat_r;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_r = shared_dat_r;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_ack = (shared_ack & (grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_ack = (shared_ack & (grant == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_err = (shared_err & (grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_err = (shared_err & (grant == 1'd1));
assign request = {(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cyc & (~monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_ack)), (monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cyc & (~monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_ack))};

// synthesis translate_off
reg dummy_d_72;
// synthesis translate_on
always @(*) begin
	slave_sel <= 5'd0;
	slave_sel[0] <= ((1'd1 & (~shared_adr[27])) & shared_adr[28]);
	slave_sel[1] <= ((1'd1 & shared_adr[27]) & shared_adr[28]);
	slave_sel[2] <= (((1'd1 & (~shared_adr[26])) & (~shared_adr[28])) & shared_adr[27]);
	slave_sel[3] <= (((1'd1 & (~shared_adr[28])) & shared_adr[26]) & shared_adr[27]);
	slave_sel[4] <= ((1'd1 & (~shared_adr[27])) & (~shared_adr[28]));
// synthesis translate_off
	dummy_d_72 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_adr = shared_adr;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_w = shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_sel = shared_sel;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_stb = shared_stb;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_we = shared_we;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cti = shared_cti;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_bte = shared_bte;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_adr = shared_adr;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_w = shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_sel = shared_sel;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_stb = shared_stb;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_we = shared_we;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_cti = shared_cti;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_bte = shared_bte;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr = shared_adr;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w = shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_sel = shared_sel;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb = shared_stb;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we = shared_we;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cti = shared_cti;
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_bte = shared_bte;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr = shared_adr;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w = shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_sel = shared_sel;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb = shared_stb;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we = shared_we;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cti = shared_cti;
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_bte = shared_bte;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_adr = shared_adr;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_w = shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_sel = shared_sel;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_stb = shared_stb;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_we = shared_we;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cti = shared_cti;
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_bte = shared_bte;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cyc = (shared_cyc & slave_sel[0]);
assign monroe_ionphoton_monroe_ionphoton_mailbox_i2_cyc = (shared_cyc & slave_sel[1]);
assign monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc = (shared_cyc & slave_sel[2]);
assign monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc = (shared_cyc & slave_sel[3]);
assign monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cyc = (shared_cyc & slave_sel[4]);
assign shared_ack = ((((monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_ack | monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack) | monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack) | monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack) | monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack);
assign shared_err = ((((monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_err | monroe_ionphoton_monroe_ionphoton_mailbox_i2_err) | monroe_ionphoton_monroe_ionphoton_csrbank0_bus_err) | monroe_ionphoton_monroe_ionphoton_csrbank1_bus_err) | monroe_ionphoton_monroe_ionphoton_csrbank2_bus_err);
assign shared_dat_r = ((((({32{slave_sel_r[0]}} & monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_r) | ({32{slave_sel_r[1]}} & monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_r)) | ({32{slave_sel_r[2]}} & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r)) | ({32{slave_sel_r[3]}} & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r)) | ({32{slave_sel_r[4]}} & monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_r));
assign monroe_ionphoton_add_identifier_adr = monroe_ionphoton_add_identifier_storage;
assign monroe_ionphoton_add_identifier_status = monroe_ionphoton_add_identifier_dat_r;
assign {user_led} = monroe_ionphoton_leds_storage;
assign monroe_ionphoton_i2c_tstriple0_o = monroe_ionphoton_i2c_out_storage[0];
assign monroe_ionphoton_i2c_tstriple0_oe = monroe_ionphoton_i2c_oe_storage[0];

// synthesis translate_off
reg dummy_d_73;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_i2c_status0 <= 2'd0;
	monroe_ionphoton_i2c_status0[0] <= monroe_ionphoton_i2c_status1;
	monroe_ionphoton_i2c_status0[1] <= monroe_ionphoton_i2c_status2;
// synthesis translate_off
	dummy_d_73 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_i2c_tstriple1_o = monroe_ionphoton_i2c_out_storage[1];
assign monroe_ionphoton_i2c_tstriple1_oe = monroe_ionphoton_i2c_oe_storage[1];
assign inout_8x0_inout_8x0_input_state = inout_8x0_serdes_i0[7];
assign inout_8x0_inout_8x0_i = (inout_8x0_serdes_i0 ^ {8{inout_8x0_inout_8x0_i_d}});
assign inout_8x0_serdes_i0 = inout_8x0_serdes_i1;
assign inout_8x0_serdes_t_in = (~inout_8x0_serdes_oe);
assign inout_8x0_serdes_o1 = inout_8x0_serdes_o0;
assign inout_8x0_serdes_pad_i1 = inout_8x0_serdes_pad_i0;
assign inout_8x0_serdes_pad_o0 = inout_8x0_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_74;
// synthesis translate_on
always @(*) begin
	inout_8x0_inout_8x0_o <= 3'd0;
	if (inout_8x0_inout_8x0_i[7]) begin
		inout_8x0_inout_8x0_o <= 3'd7;
	end
	if (inout_8x0_inout_8x0_i[6]) begin
		inout_8x0_inout_8x0_o <= 3'd6;
	end
	if (inout_8x0_inout_8x0_i[5]) begin
		inout_8x0_inout_8x0_o <= 3'd5;
	end
	if (inout_8x0_inout_8x0_i[4]) begin
		inout_8x0_inout_8x0_o <= 3'd4;
	end
	if (inout_8x0_inout_8x0_i[3]) begin
		inout_8x0_inout_8x0_o <= 2'd3;
	end
	if (inout_8x0_inout_8x0_i[2]) begin
		inout_8x0_inout_8x0_o <= 2'd2;
	end
	if (inout_8x0_inout_8x0_i[1]) begin
		inout_8x0_inout_8x0_o <= 1'd1;
	end
	if (inout_8x0_inout_8x0_i[0]) begin
		inout_8x0_inout_8x0_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_74 <= dummy_s;
// synthesis translate_on
end
assign inout_8x0_inout_8x0_n = (inout_8x0_inout_8x0_i == 1'd0);
assign inout_8x1_inout_8x1_input_state = inout_8x1_serdes_i0[7];
assign inout_8x1_inout_8x1_i = (inout_8x1_serdes_i0 ^ {8{inout_8x1_inout_8x1_i_d}});
assign inout_8x1_serdes_i0 = inout_8x1_serdes_i1;
assign inout_8x1_serdes_t_in = (~inout_8x1_serdes_oe);
assign inout_8x1_serdes_o1 = inout_8x1_serdes_o0;
assign inout_8x1_serdes_pad_i1 = inout_8x1_serdes_pad_i0;
assign inout_8x1_serdes_pad_o0 = inout_8x1_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_75;
// synthesis translate_on
always @(*) begin
	inout_8x1_inout_8x1_o <= 3'd0;
	if (inout_8x1_inout_8x1_i[7]) begin
		inout_8x1_inout_8x1_o <= 3'd7;
	end
	if (inout_8x1_inout_8x1_i[6]) begin
		inout_8x1_inout_8x1_o <= 3'd6;
	end
	if (inout_8x1_inout_8x1_i[5]) begin
		inout_8x1_inout_8x1_o <= 3'd5;
	end
	if (inout_8x1_inout_8x1_i[4]) begin
		inout_8x1_inout_8x1_o <= 3'd4;
	end
	if (inout_8x1_inout_8x1_i[3]) begin
		inout_8x1_inout_8x1_o <= 2'd3;
	end
	if (inout_8x1_inout_8x1_i[2]) begin
		inout_8x1_inout_8x1_o <= 2'd2;
	end
	if (inout_8x1_inout_8x1_i[1]) begin
		inout_8x1_inout_8x1_o <= 1'd1;
	end
	if (inout_8x1_inout_8x1_i[0]) begin
		inout_8x1_inout_8x1_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_75 <= dummy_s;
// synthesis translate_on
end
assign inout_8x1_inout_8x1_n = (inout_8x1_inout_8x1_i == 1'd0);
assign inout_8x2_inout_8x2_input_state = inout_8x2_serdes_i0[7];
assign inout_8x2_inout_8x2_i = (inout_8x2_serdes_i0 ^ {8{inout_8x2_inout_8x2_i_d}});
assign inout_8x2_serdes_i0 = inout_8x2_serdes_i1;
assign inout_8x2_serdes_t_in = (~inout_8x2_serdes_oe);
assign inout_8x2_serdes_o1 = inout_8x2_serdes_o0;
assign inout_8x2_serdes_pad_i1 = inout_8x2_serdes_pad_i0;
assign inout_8x2_serdes_pad_o0 = inout_8x2_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_76;
// synthesis translate_on
always @(*) begin
	inout_8x2_inout_8x2_o <= 3'd0;
	if (inout_8x2_inout_8x2_i[7]) begin
		inout_8x2_inout_8x2_o <= 3'd7;
	end
	if (inout_8x2_inout_8x2_i[6]) begin
		inout_8x2_inout_8x2_o <= 3'd6;
	end
	if (inout_8x2_inout_8x2_i[5]) begin
		inout_8x2_inout_8x2_o <= 3'd5;
	end
	if (inout_8x2_inout_8x2_i[4]) begin
		inout_8x2_inout_8x2_o <= 3'd4;
	end
	if (inout_8x2_inout_8x2_i[3]) begin
		inout_8x2_inout_8x2_o <= 2'd3;
	end
	if (inout_8x2_inout_8x2_i[2]) begin
		inout_8x2_inout_8x2_o <= 2'd2;
	end
	if (inout_8x2_inout_8x2_i[1]) begin
		inout_8x2_inout_8x2_o <= 1'd1;
	end
	if (inout_8x2_inout_8x2_i[0]) begin
		inout_8x2_inout_8x2_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_76 <= dummy_s;
// synthesis translate_on
end
assign inout_8x2_inout_8x2_n = (inout_8x2_inout_8x2_i == 1'd0);
assign inout_8x3_inout_8x3_input_state = inout_8x3_serdes_i0[7];
assign inout_8x3_inout_8x3_i = (inout_8x3_serdes_i0 ^ {8{inout_8x3_inout_8x3_i_d}});
assign inout_8x3_serdes_i0 = inout_8x3_serdes_i1;
assign inout_8x3_serdes_t_in = (~inout_8x3_serdes_oe);
assign inout_8x3_serdes_o1 = inout_8x3_serdes_o0;
assign inout_8x3_serdes_pad_i1 = inout_8x3_serdes_pad_i0;
assign inout_8x3_serdes_pad_o0 = inout_8x3_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_77;
// synthesis translate_on
always @(*) begin
	inout_8x3_inout_8x3_o <= 3'd0;
	if (inout_8x3_inout_8x3_i[7]) begin
		inout_8x3_inout_8x3_o <= 3'd7;
	end
	if (inout_8x3_inout_8x3_i[6]) begin
		inout_8x3_inout_8x3_o <= 3'd6;
	end
	if (inout_8x3_inout_8x3_i[5]) begin
		inout_8x3_inout_8x3_o <= 3'd5;
	end
	if (inout_8x3_inout_8x3_i[4]) begin
		inout_8x3_inout_8x3_o <= 3'd4;
	end
	if (inout_8x3_inout_8x3_i[3]) begin
		inout_8x3_inout_8x3_o <= 2'd3;
	end
	if (inout_8x3_inout_8x3_i[2]) begin
		inout_8x3_inout_8x3_o <= 2'd2;
	end
	if (inout_8x3_inout_8x3_i[1]) begin
		inout_8x3_inout_8x3_o <= 1'd1;
	end
	if (inout_8x3_inout_8x3_i[0]) begin
		inout_8x3_inout_8x3_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_77 <= dummy_s;
// synthesis translate_on
end
assign inout_8x3_inout_8x3_n = (inout_8x3_inout_8x3_i == 1'd0);
assign spimaster0_spimachine0_length = spimaster0_config_length;
assign spimaster0_spimachine0_end0 = spimaster0_config_end;
assign spimaster0_spimachine0_div = spimaster0_config_div;
assign spimaster0_spimachine0_clk_phase = spimaster0_config_clk_phase;
assign spimaster0_spimachine0_lsb_first = spimaster0_config_lsb_first;
assign spimaster0_interface_half_duplex = spimaster0_config_half_duplex;
assign spimaster0_interface_cs0 = spimaster0_config_cs;
assign spimaster0_interface_cs_polarity = {3{spimaster0_config_cs_polarity}};
assign spimaster0_interface_clk_polarity = spimaster0_config_clk_polarity;
assign spimaster0_interface_offline = spimaster0_config_offline;
assign spimaster0_interface_cs_next = spimaster0_spimachine0_cs_next;
assign spimaster0_interface_clk_next = spimaster0_spimachine0_clk_next;
assign spimaster0_interface_ce = spimaster0_spimachine0_ce;
assign spimaster0_interface_sample = spimaster0_spimachine0_sample;
assign spimaster0_spimachine0_sdi = spimaster0_interface_sdi;
assign spimaster0_interface_sdo = spimaster0_spimachine0_sdo;
assign spimaster0_spimachine0_load0 = ((spimaster0_ointerface0_stb & spimaster0_spimachine0_writable) & (~spimaster0_ointerface0_address));
assign spimaster0_spimachine0_pdo = spimaster0_ointerface0_data;
assign spimaster0_ointerface0_busy = (~spimaster0_spimachine0_writable);
assign spimaster0_iinterface0_stb = (spimaster0_spimachine0_readable & spimaster0_read);
assign spimaster0_iinterface0_data = spimaster0_spimachine0_pdi;
assign spimaster0_interface_sdi = (spimaster0_interface_half_duplex ? spimaster0_interface_mosi_reg : spimaster0_interface_miso_reg);
assign spimaster0_spimachine0_ce = (spimaster0_spimachine0_done & spimaster0_spimachine0_count);
assign spimaster0_spimachine0_pdi = (spimaster0_spimachine0_lsb_first ? {spimaster0_spimachine0_sdi, spimaster0_spimachine0_sr[31:1]} : {spimaster0_spimachine0_sr[30:0], spimaster0_spimachine0_sdi});
assign spimaster0_spimachine0_cnt_done = (spimaster0_spimachine0_cnt == 1'd0);
assign spimaster0_spimachine0_done = (spimaster0_spimachine0_cnt_done & (~spimaster0_spimachine0_do_extend));

// synthesis translate_off
reg dummy_d_78;
// synthesis translate_on
always @(*) begin
	spimaster0_spimachine0_clk_next <= 1'd0;
	spimaster0_spimachine0_cs_next <= 1'd0;
	spimaster0_spimachine0_idle <= 1'd0;
	spimaster0_spimachine0_readable <= 1'd0;
	spimaster0_spimachine0_writable <= 1'd0;
	spimaster0_spimachine0_load1 <= 1'd0;
	spimaster0_spimachine0_shift <= 1'd0;
	spimaster0_spimachine0_sample <= 1'd0;
	spimaster0_spimachine0_extend <= 1'd0;
	spimaster0_spimachine0_count <= 1'd0;
	spimaster0_next_state <= 3'd0;
	spimaster0_next_state <= spimaster0_state;
	case (spimaster0_state)
		1'd1: begin
			spimaster0_spimachine0_cs_next <= 1'd1;
			spimaster0_spimachine0_count <= 1'd1;
			spimaster0_spimachine0_extend <= 1'd1;
			spimaster0_spimachine0_clk_next <= 1'd1;
			if (spimaster0_spimachine0_done) begin
				spimaster0_next_state <= 2'd2;
			end
		end
		2'd2: begin
			spimaster0_spimachine0_cs_next <= 1'd1;
			spimaster0_spimachine0_count <= 1'd1;
			spimaster0_spimachine0_clk_next <= (~spimaster0_spimachine0_clk_phase);
			if (spimaster0_spimachine0_done) begin
				spimaster0_spimachine0_sample <= 1'd1;
				spimaster0_next_state <= 2'd3;
			end
		end
		2'd3: begin
			spimaster0_spimachine0_cs_next <= 1'd1;
			spimaster0_spimachine0_count <= 1'd1;
			spimaster0_spimachine0_extend <= 1'd1;
			spimaster0_spimachine0_clk_next <= spimaster0_spimachine0_clk_phase;
			if (spimaster0_spimachine0_done) begin
				if ((spimaster0_spimachine0_n == 1'd0)) begin
					spimaster0_spimachine0_readable <= 1'd1;
					spimaster0_spimachine0_writable <= 1'd1;
					if (spimaster0_spimachine0_end1) begin
						spimaster0_spimachine0_clk_next <= 1'd0;
						spimaster0_spimachine0_writable <= 1'd0;
						if (spimaster0_spimachine0_clk_phase) begin
							spimaster0_spimachine0_cs_next <= 1'd0;
							spimaster0_next_state <= 3'd5;
						end else begin
							spimaster0_next_state <= 3'd4;
						end
					end else begin
						if (spimaster0_spimachine0_load0) begin
							spimaster0_spimachine0_load1 <= 1'd1;
							spimaster0_next_state <= 2'd2;
						end else begin
							spimaster0_spimachine0_count <= 1'd0;
						end
					end
				end else begin
					spimaster0_spimachine0_shift <= 1'd1;
					spimaster0_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			spimaster0_spimachine0_count <= 1'd1;
			if (spimaster0_spimachine0_done) begin
				spimaster0_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (spimaster0_spimachine0_done) begin
				spimaster0_next_state <= 1'd0;
			end else begin
				spimaster0_spimachine0_count <= 1'd1;
			end
		end
		default: begin
			spimaster0_spimachine0_idle <= 1'd1;
			spimaster0_spimachine0_writable <= 1'd1;
			spimaster0_spimachine0_cs_next <= 1'd1;
			if (spimaster0_spimachine0_load0) begin
				spimaster0_spimachine0_count <= 1'd1;
				spimaster0_spimachine0_load1 <= 1'd1;
				if (spimaster0_spimachine0_clk_phase) begin
					spimaster0_next_state <= 1'd1;
				end else begin
					spimaster0_spimachine0_extend <= 1'd1;
					spimaster0_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_78 <= dummy_s;
// synthesis translate_on
end
assign spimaster1_spimachine1_length = spimaster1_config_length;
assign spimaster1_spimachine1_end0 = spimaster1_config_end;
assign spimaster1_spimachine1_div = spimaster1_config_div;
assign spimaster1_spimachine1_clk_phase = spimaster1_config_clk_phase;
assign spimaster1_spimachine1_lsb_first = spimaster1_config_lsb_first;
assign spimaster1_interface_half_duplex = spimaster1_config_half_duplex;
assign spimaster1_interface_cs0 = spimaster1_config_cs;
assign spimaster1_interface_cs_polarity = {3{spimaster1_config_cs_polarity}};
assign spimaster1_interface_clk_polarity = spimaster1_config_clk_polarity;
assign spimaster1_interface_offline = spimaster1_config_offline;
assign spimaster1_interface_cs_next = spimaster1_spimachine1_cs_next;
assign spimaster1_interface_clk_next = spimaster1_spimachine1_clk_next;
assign spimaster1_interface_ce = spimaster1_spimachine1_ce;
assign spimaster1_interface_sample = spimaster1_spimachine1_sample;
assign spimaster1_spimachine1_sdi = spimaster1_interface_sdi;
assign spimaster1_interface_sdo = spimaster1_spimachine1_sdo;
assign spimaster1_spimachine1_load0 = ((spimaster1_ointerface1_stb & spimaster1_spimachine1_writable) & (~spimaster1_ointerface1_address));
assign spimaster1_spimachine1_pdo = spimaster1_ointerface1_data;
assign spimaster1_ointerface1_busy = (~spimaster1_spimachine1_writable);
assign spimaster1_iinterface1_stb = (spimaster1_spimachine1_readable & spimaster1_read);
assign spimaster1_iinterface1_data = spimaster1_spimachine1_pdi;
assign spimaster1_interface_sdi = (spimaster1_interface_half_duplex ? spimaster1_interface_mosi_reg : spimaster1_interface_miso_reg);
assign spimaster1_spimachine1_ce = (spimaster1_spimachine1_done & spimaster1_spimachine1_count);
assign spimaster1_spimachine1_pdi = (spimaster1_spimachine1_lsb_first ? {spimaster1_spimachine1_sdi, spimaster1_spimachine1_sr[31:1]} : {spimaster1_spimachine1_sr[30:0], spimaster1_spimachine1_sdi});
assign spimaster1_spimachine1_cnt_done = (spimaster1_spimachine1_cnt == 1'd0);
assign spimaster1_spimachine1_done = (spimaster1_spimachine1_cnt_done & (~spimaster1_spimachine1_do_extend));

// synthesis translate_off
reg dummy_d_79;
// synthesis translate_on
always @(*) begin
	spimaster1_spimachine1_clk_next <= 1'd0;
	spimaster1_spimachine1_cs_next <= 1'd0;
	spimaster1_spimachine1_idle <= 1'd0;
	spimaster1_spimachine1_readable <= 1'd0;
	spimaster1_spimachine1_writable <= 1'd0;
	spimaster1_spimachine1_load1 <= 1'd0;
	spimaster1_spimachine1_shift <= 1'd0;
	spimaster1_spimachine1_sample <= 1'd0;
	spimaster1_spimachine1_extend <= 1'd0;
	spimaster1_spimachine1_count <= 1'd0;
	spimaster1_next_state <= 3'd0;
	spimaster1_next_state <= spimaster1_state;
	case (spimaster1_state)
		1'd1: begin
			spimaster1_spimachine1_cs_next <= 1'd1;
			spimaster1_spimachine1_count <= 1'd1;
			spimaster1_spimachine1_extend <= 1'd1;
			spimaster1_spimachine1_clk_next <= 1'd1;
			if (spimaster1_spimachine1_done) begin
				spimaster1_next_state <= 2'd2;
			end
		end
		2'd2: begin
			spimaster1_spimachine1_cs_next <= 1'd1;
			spimaster1_spimachine1_count <= 1'd1;
			spimaster1_spimachine1_clk_next <= (~spimaster1_spimachine1_clk_phase);
			if (spimaster1_spimachine1_done) begin
				spimaster1_spimachine1_sample <= 1'd1;
				spimaster1_next_state <= 2'd3;
			end
		end
		2'd3: begin
			spimaster1_spimachine1_cs_next <= 1'd1;
			spimaster1_spimachine1_count <= 1'd1;
			spimaster1_spimachine1_extend <= 1'd1;
			spimaster1_spimachine1_clk_next <= spimaster1_spimachine1_clk_phase;
			if (spimaster1_spimachine1_done) begin
				if ((spimaster1_spimachine1_n == 1'd0)) begin
					spimaster1_spimachine1_readable <= 1'd1;
					spimaster1_spimachine1_writable <= 1'd1;
					if (spimaster1_spimachine1_end1) begin
						spimaster1_spimachine1_clk_next <= 1'd0;
						spimaster1_spimachine1_writable <= 1'd0;
						if (spimaster1_spimachine1_clk_phase) begin
							spimaster1_spimachine1_cs_next <= 1'd0;
							spimaster1_next_state <= 3'd5;
						end else begin
							spimaster1_next_state <= 3'd4;
						end
					end else begin
						if (spimaster1_spimachine1_load0) begin
							spimaster1_spimachine1_load1 <= 1'd1;
							spimaster1_next_state <= 2'd2;
						end else begin
							spimaster1_spimachine1_count <= 1'd0;
						end
					end
				end else begin
					spimaster1_spimachine1_shift <= 1'd1;
					spimaster1_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			spimaster1_spimachine1_count <= 1'd1;
			if (spimaster1_spimachine1_done) begin
				spimaster1_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (spimaster1_spimachine1_done) begin
				spimaster1_next_state <= 1'd0;
			end else begin
				spimaster1_spimachine1_count <= 1'd1;
			end
		end
		default: begin
			spimaster1_spimachine1_idle <= 1'd1;
			spimaster1_spimachine1_writable <= 1'd1;
			spimaster1_spimachine1_cs_next <= 1'd1;
			if (spimaster1_spimachine1_load0) begin
				spimaster1_spimachine1_count <= 1'd1;
				spimaster1_spimachine1_load1 <= 1'd1;
				if (spimaster1_spimachine1_clk_phase) begin
					spimaster1_next_state <= 1'd1;
				end else begin
					spimaster1_spimachine1_extend <= 1'd1;
					spimaster1_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_79 <= dummy_s;
// synthesis translate_on
end
assign spimaster2_spimachine2_length = spimaster2_config_length;
assign spimaster2_spimachine2_end0 = spimaster2_config_end;
assign spimaster2_spimachine2_div = spimaster2_config_div;
assign spimaster2_spimachine2_clk_phase = spimaster2_config_clk_phase;
assign spimaster2_spimachine2_lsb_first = spimaster2_config_lsb_first;
assign spimaster2_interface_half_duplex = spimaster2_config_half_duplex;
assign spimaster2_interface_cs0 = spimaster2_config_cs;
assign spimaster2_interface_cs_polarity = {3{spimaster2_config_cs_polarity}};
assign spimaster2_interface_clk_polarity = spimaster2_config_clk_polarity;
assign spimaster2_interface_offline = spimaster2_config_offline;
assign spimaster2_interface_cs_next = spimaster2_spimachine2_cs_next;
assign spimaster2_interface_clk_next = spimaster2_spimachine2_clk_next;
assign spimaster2_interface_ce = spimaster2_spimachine2_ce;
assign spimaster2_interface_sample = spimaster2_spimachine2_sample;
assign spimaster2_spimachine2_sdi = spimaster2_interface_sdi;
assign spimaster2_interface_sdo = spimaster2_spimachine2_sdo;
assign spimaster2_spimachine2_load0 = ((spimaster2_ointerface2_stb & spimaster2_spimachine2_writable) & (~spimaster2_ointerface2_address));
assign spimaster2_spimachine2_pdo = spimaster2_ointerface2_data;
assign spimaster2_ointerface2_busy = (~spimaster2_spimachine2_writable);
assign spimaster2_iinterface2_stb = (spimaster2_spimachine2_readable & spimaster2_read);
assign spimaster2_iinterface2_data = spimaster2_spimachine2_pdi;
assign spimaster2_interface_sdi = (spimaster2_interface_half_duplex ? spimaster2_interface_mosi_reg : spimaster2_interface_miso_reg);
assign spimaster2_spimachine2_ce = (spimaster2_spimachine2_done & spimaster2_spimachine2_count);
assign spimaster2_spimachine2_pdi = (spimaster2_spimachine2_lsb_first ? {spimaster2_spimachine2_sdi, spimaster2_spimachine2_sr[31:1]} : {spimaster2_spimachine2_sr[30:0], spimaster2_spimachine2_sdi});
assign spimaster2_spimachine2_cnt_done = (spimaster2_spimachine2_cnt == 1'd0);
assign spimaster2_spimachine2_done = (spimaster2_spimachine2_cnt_done & (~spimaster2_spimachine2_do_extend));

// synthesis translate_off
reg dummy_d_80;
// synthesis translate_on
always @(*) begin
	spimaster2_spimachine2_clk_next <= 1'd0;
	spimaster2_spimachine2_cs_next <= 1'd0;
	spimaster2_spimachine2_idle <= 1'd0;
	spimaster2_spimachine2_readable <= 1'd0;
	spimaster2_spimachine2_writable <= 1'd0;
	spimaster2_spimachine2_load1 <= 1'd0;
	spimaster2_spimachine2_shift <= 1'd0;
	spimaster2_spimachine2_sample <= 1'd0;
	spimaster2_spimachine2_extend <= 1'd0;
	spimaster2_spimachine2_count <= 1'd0;
	spimaster2_next_state <= 3'd0;
	spimaster2_next_state <= spimaster2_state;
	case (spimaster2_state)
		1'd1: begin
			spimaster2_spimachine2_cs_next <= 1'd1;
			spimaster2_spimachine2_count <= 1'd1;
			spimaster2_spimachine2_extend <= 1'd1;
			spimaster2_spimachine2_clk_next <= 1'd1;
			if (spimaster2_spimachine2_done) begin
				spimaster2_next_state <= 2'd2;
			end
		end
		2'd2: begin
			spimaster2_spimachine2_cs_next <= 1'd1;
			spimaster2_spimachine2_count <= 1'd1;
			spimaster2_spimachine2_clk_next <= (~spimaster2_spimachine2_clk_phase);
			if (spimaster2_spimachine2_done) begin
				spimaster2_spimachine2_sample <= 1'd1;
				spimaster2_next_state <= 2'd3;
			end
		end
		2'd3: begin
			spimaster2_spimachine2_cs_next <= 1'd1;
			spimaster2_spimachine2_count <= 1'd1;
			spimaster2_spimachine2_extend <= 1'd1;
			spimaster2_spimachine2_clk_next <= spimaster2_spimachine2_clk_phase;
			if (spimaster2_spimachine2_done) begin
				if ((spimaster2_spimachine2_n == 1'd0)) begin
					spimaster2_spimachine2_readable <= 1'd1;
					spimaster2_spimachine2_writable <= 1'd1;
					if (spimaster2_spimachine2_end1) begin
						spimaster2_spimachine2_clk_next <= 1'd0;
						spimaster2_spimachine2_writable <= 1'd0;
						if (spimaster2_spimachine2_clk_phase) begin
							spimaster2_spimachine2_cs_next <= 1'd0;
							spimaster2_next_state <= 3'd5;
						end else begin
							spimaster2_next_state <= 3'd4;
						end
					end else begin
						if (spimaster2_spimachine2_load0) begin
							spimaster2_spimachine2_load1 <= 1'd1;
							spimaster2_next_state <= 2'd2;
						end else begin
							spimaster2_spimachine2_count <= 1'd0;
						end
					end
				end else begin
					spimaster2_spimachine2_shift <= 1'd1;
					spimaster2_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			spimaster2_spimachine2_count <= 1'd1;
			if (spimaster2_spimachine2_done) begin
				spimaster2_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (spimaster2_spimachine2_done) begin
				spimaster2_next_state <= 1'd0;
			end else begin
				spimaster2_spimachine2_count <= 1'd1;
			end
		end
		default: begin
			spimaster2_spimachine2_idle <= 1'd1;
			spimaster2_spimachine2_writable <= 1'd1;
			spimaster2_spimachine2_cs_next <= 1'd1;
			if (spimaster2_spimachine2_load0) begin
				spimaster2_spimachine2_count <= 1'd1;
				spimaster2_spimachine2_load1 <= 1'd1;
				if (spimaster2_spimachine2_clk_phase) begin
					spimaster2_next_state <= 1'd1;
				end else begin
					spimaster2_spimachine2_extend <= 1'd1;
					spimaster2_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_80 <= dummy_s;
// synthesis translate_on
end
assign sfp_ctl_led_1 = output0_pad_o;
assign sfp_ctl_led_2 = output1_pad_o;
assign monroe_ionphoton_rtio_tsc_i = monroe_ionphoton_rtio_tsc_coarse_ts;
assign monroe_ionphoton_rtio_tsc_coarse_ts_sys = monroe_ionphoton_rtio_tsc_o;
assign monroe_ionphoton_rtio_tsc_full_ts = (monroe_ionphoton_rtio_tsc_coarse_ts <<< 2'd3);
assign monroe_ionphoton_rtio_tsc_full_ts_sys = (monroe_ionphoton_rtio_tsc_coarse_ts_sys <<< 2'd3);

// synthesis translate_off
reg dummy_d_81;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_tsc_value_sys <= 61'd0;
	monroe_ionphoton_rtio_tsc_value_sys[60] <= monroe_ionphoton_rtio_tsc_value_gray_sys[60];
	monroe_ionphoton_rtio_tsc_value_sys[59] <= (monroe_ionphoton_rtio_tsc_value_sys[60] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[59]);
	monroe_ionphoton_rtio_tsc_value_sys[58] <= (monroe_ionphoton_rtio_tsc_value_sys[59] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[58]);
	monroe_ionphoton_rtio_tsc_value_sys[57] <= (monroe_ionphoton_rtio_tsc_value_sys[58] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[57]);
	monroe_ionphoton_rtio_tsc_value_sys[56] <= (monroe_ionphoton_rtio_tsc_value_sys[57] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[56]);
	monroe_ionphoton_rtio_tsc_value_sys[55] <= (monroe_ionphoton_rtio_tsc_value_sys[56] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[55]);
	monroe_ionphoton_rtio_tsc_value_sys[54] <= (monroe_ionphoton_rtio_tsc_value_sys[55] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[54]);
	monroe_ionphoton_rtio_tsc_value_sys[53] <= (monroe_ionphoton_rtio_tsc_value_sys[54] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[53]);
	monroe_ionphoton_rtio_tsc_value_sys[52] <= (monroe_ionphoton_rtio_tsc_value_sys[53] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[52]);
	monroe_ionphoton_rtio_tsc_value_sys[51] <= (monroe_ionphoton_rtio_tsc_value_sys[52] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[51]);
	monroe_ionphoton_rtio_tsc_value_sys[50] <= (monroe_ionphoton_rtio_tsc_value_sys[51] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[50]);
	monroe_ionphoton_rtio_tsc_value_sys[49] <= (monroe_ionphoton_rtio_tsc_value_sys[50] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[49]);
	monroe_ionphoton_rtio_tsc_value_sys[48] <= (monroe_ionphoton_rtio_tsc_value_sys[49] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[48]);
	monroe_ionphoton_rtio_tsc_value_sys[47] <= (monroe_ionphoton_rtio_tsc_value_sys[48] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[47]);
	monroe_ionphoton_rtio_tsc_value_sys[46] <= (monroe_ionphoton_rtio_tsc_value_sys[47] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[46]);
	monroe_ionphoton_rtio_tsc_value_sys[45] <= (monroe_ionphoton_rtio_tsc_value_sys[46] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[45]);
	monroe_ionphoton_rtio_tsc_value_sys[44] <= (monroe_ionphoton_rtio_tsc_value_sys[45] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[44]);
	monroe_ionphoton_rtio_tsc_value_sys[43] <= (monroe_ionphoton_rtio_tsc_value_sys[44] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[43]);
	monroe_ionphoton_rtio_tsc_value_sys[42] <= (monroe_ionphoton_rtio_tsc_value_sys[43] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[42]);
	monroe_ionphoton_rtio_tsc_value_sys[41] <= (monroe_ionphoton_rtio_tsc_value_sys[42] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[41]);
	monroe_ionphoton_rtio_tsc_value_sys[40] <= (monroe_ionphoton_rtio_tsc_value_sys[41] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[40]);
	monroe_ionphoton_rtio_tsc_value_sys[39] <= (monroe_ionphoton_rtio_tsc_value_sys[40] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[39]);
	monroe_ionphoton_rtio_tsc_value_sys[38] <= (monroe_ionphoton_rtio_tsc_value_sys[39] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[38]);
	monroe_ionphoton_rtio_tsc_value_sys[37] <= (monroe_ionphoton_rtio_tsc_value_sys[38] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[37]);
	monroe_ionphoton_rtio_tsc_value_sys[36] <= (monroe_ionphoton_rtio_tsc_value_sys[37] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[36]);
	monroe_ionphoton_rtio_tsc_value_sys[35] <= (monroe_ionphoton_rtio_tsc_value_sys[36] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[35]);
	monroe_ionphoton_rtio_tsc_value_sys[34] <= (monroe_ionphoton_rtio_tsc_value_sys[35] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[34]);
	monroe_ionphoton_rtio_tsc_value_sys[33] <= (monroe_ionphoton_rtio_tsc_value_sys[34] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[33]);
	monroe_ionphoton_rtio_tsc_value_sys[32] <= (monroe_ionphoton_rtio_tsc_value_sys[33] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[32]);
	monroe_ionphoton_rtio_tsc_value_sys[31] <= (monroe_ionphoton_rtio_tsc_value_sys[32] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[31]);
	monroe_ionphoton_rtio_tsc_value_sys[30] <= (monroe_ionphoton_rtio_tsc_value_sys[31] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[30]);
	monroe_ionphoton_rtio_tsc_value_sys[29] <= (monroe_ionphoton_rtio_tsc_value_sys[30] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[29]);
	monroe_ionphoton_rtio_tsc_value_sys[28] <= (monroe_ionphoton_rtio_tsc_value_sys[29] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[28]);
	monroe_ionphoton_rtio_tsc_value_sys[27] <= (monroe_ionphoton_rtio_tsc_value_sys[28] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[27]);
	monroe_ionphoton_rtio_tsc_value_sys[26] <= (monroe_ionphoton_rtio_tsc_value_sys[27] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[26]);
	monroe_ionphoton_rtio_tsc_value_sys[25] <= (monroe_ionphoton_rtio_tsc_value_sys[26] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[25]);
	monroe_ionphoton_rtio_tsc_value_sys[24] <= (monroe_ionphoton_rtio_tsc_value_sys[25] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[24]);
	monroe_ionphoton_rtio_tsc_value_sys[23] <= (monroe_ionphoton_rtio_tsc_value_sys[24] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[23]);
	monroe_ionphoton_rtio_tsc_value_sys[22] <= (monroe_ionphoton_rtio_tsc_value_sys[23] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[22]);
	monroe_ionphoton_rtio_tsc_value_sys[21] <= (monroe_ionphoton_rtio_tsc_value_sys[22] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[21]);
	monroe_ionphoton_rtio_tsc_value_sys[20] <= (monroe_ionphoton_rtio_tsc_value_sys[21] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[20]);
	monroe_ionphoton_rtio_tsc_value_sys[19] <= (monroe_ionphoton_rtio_tsc_value_sys[20] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[19]);
	monroe_ionphoton_rtio_tsc_value_sys[18] <= (monroe_ionphoton_rtio_tsc_value_sys[19] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[18]);
	monroe_ionphoton_rtio_tsc_value_sys[17] <= (monroe_ionphoton_rtio_tsc_value_sys[18] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[17]);
	monroe_ionphoton_rtio_tsc_value_sys[16] <= (monroe_ionphoton_rtio_tsc_value_sys[17] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[16]);
	monroe_ionphoton_rtio_tsc_value_sys[15] <= (monroe_ionphoton_rtio_tsc_value_sys[16] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[15]);
	monroe_ionphoton_rtio_tsc_value_sys[14] <= (monroe_ionphoton_rtio_tsc_value_sys[15] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[14]);
	monroe_ionphoton_rtio_tsc_value_sys[13] <= (monroe_ionphoton_rtio_tsc_value_sys[14] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[13]);
	monroe_ionphoton_rtio_tsc_value_sys[12] <= (monroe_ionphoton_rtio_tsc_value_sys[13] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[12]);
	monroe_ionphoton_rtio_tsc_value_sys[11] <= (monroe_ionphoton_rtio_tsc_value_sys[12] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[11]);
	monroe_ionphoton_rtio_tsc_value_sys[10] <= (monroe_ionphoton_rtio_tsc_value_sys[11] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[10]);
	monroe_ionphoton_rtio_tsc_value_sys[9] <= (monroe_ionphoton_rtio_tsc_value_sys[10] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[9]);
	monroe_ionphoton_rtio_tsc_value_sys[8] <= (monroe_ionphoton_rtio_tsc_value_sys[9] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[8]);
	monroe_ionphoton_rtio_tsc_value_sys[7] <= (monroe_ionphoton_rtio_tsc_value_sys[8] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[7]);
	monroe_ionphoton_rtio_tsc_value_sys[6] <= (monroe_ionphoton_rtio_tsc_value_sys[7] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[6]);
	monroe_ionphoton_rtio_tsc_value_sys[5] <= (monroe_ionphoton_rtio_tsc_value_sys[6] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[5]);
	monroe_ionphoton_rtio_tsc_value_sys[4] <= (monroe_ionphoton_rtio_tsc_value_sys[5] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[4]);
	monroe_ionphoton_rtio_tsc_value_sys[3] <= (monroe_ionphoton_rtio_tsc_value_sys[4] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[3]);
	monroe_ionphoton_rtio_tsc_value_sys[2] <= (monroe_ionphoton_rtio_tsc_value_sys[3] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[2]);
	monroe_ionphoton_rtio_tsc_value_sys[1] <= (monroe_ionphoton_rtio_tsc_value_sys[2] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[1]);
	monroe_ionphoton_rtio_tsc_value_sys[0] <= (monroe_ionphoton_rtio_tsc_value_sys[1] ^ monroe_ionphoton_rtio_tsc_value_gray_sys[0]);
// synthesis translate_off
	dummy_d_81 <= dummy_s;
// synthesis translate_on
end
assign rsys_clk = sys_clk;
assign rsys_rst = monroe_ionphoton_rtio_core_cmd_reset;
assign rio_clk = rtio_clk;
assign rio_phy_clk = rtio_clk;
assign monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp = monroe_ionphoton_rtio_tsc_coarse_ts;
assign monroe_ionphoton_rtio_core_async_error_w = {monroe_ionphoton_rtio_core_o_sequence_error, monroe_ionphoton_rtio_core_o_busy, monroe_ionphoton_rtio_core_o_collision};
assign monroe_ionphoton_rtio_core_o_collision_sync_i = monroe_ionphoton_rtio_core_outputs_collision;
assign monroe_ionphoton_rtio_core_o_collision_sync_data_i = monroe_ionphoton_rtio_core_outputs_collision_channel;
assign monroe_ionphoton_rtio_core_o_busy_sync_i = monroe_ionphoton_rtio_core_outputs_busy;
assign monroe_ionphoton_rtio_core_o_busy_sync_data_i = monroe_ionphoton_rtio_core_outputs_busy_channel;
assign monroe_ionphoton_rtio_core_outputs_record0_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_writable = monroe_ionphoton_rtio_core_outputs_record0_writable;
assign monroe_ionphoton_rtio_core_outputs_record0_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_seqn;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record1_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_writable = monroe_ionphoton_rtio_core_outputs_record1_writable;
assign monroe_ionphoton_rtio_core_outputs_record1_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_seqn;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record2_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_writable = monroe_ionphoton_rtio_core_outputs_record2_writable;
assign monroe_ionphoton_rtio_core_outputs_record2_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_seqn;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record3_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_writable = monroe_ionphoton_rtio_core_outputs_record3_writable;
assign monroe_ionphoton_rtio_core_outputs_record3_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_seqn;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record4_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_writable = monroe_ionphoton_rtio_core_outputs_record4_writable;
assign monroe_ionphoton_rtio_core_outputs_record4_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_seqn;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record5_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_writable = monroe_ionphoton_rtio_core_outputs_record5_writable;
assign monroe_ionphoton_rtio_core_outputs_record5_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_seqn;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record6_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_writable = monroe_ionphoton_rtio_core_outputs_record6_writable;
assign monroe_ionphoton_rtio_core_outputs_record6_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_seqn;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record7_we = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_we;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_writable = monroe_ionphoton_rtio_core_outputs_record7_writable;
assign monroe_ionphoton_rtio_core_outputs_record7_seqn0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_seqn;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_channel0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_address0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_address;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_data0 = monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_data;
assign monroe_ionphoton_rtio_core_outputs_record0_re = monroe_ionphoton_rtio_core_outputs_gates_record0_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_readable = monroe_ionphoton_rtio_core_outputs_record0_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_seqn0 = monroe_ionphoton_rtio_core_outputs_record0_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record0_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address0 = monroe_ionphoton_rtio_core_outputs_record0_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data0 = monroe_ionphoton_rtio_core_outputs_record0_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record1_re = monroe_ionphoton_rtio_core_outputs_gates_record1_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_readable = monroe_ionphoton_rtio_core_outputs_record1_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_seqn0 = monroe_ionphoton_rtio_core_outputs_record1_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record1_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address0 = monroe_ionphoton_rtio_core_outputs_record1_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data0 = monroe_ionphoton_rtio_core_outputs_record1_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record2_re = monroe_ionphoton_rtio_core_outputs_gates_record2_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_readable = monroe_ionphoton_rtio_core_outputs_record2_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_seqn0 = monroe_ionphoton_rtio_core_outputs_record2_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record2_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address0 = monroe_ionphoton_rtio_core_outputs_record2_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data0 = monroe_ionphoton_rtio_core_outputs_record2_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record3_re = monroe_ionphoton_rtio_core_outputs_gates_record3_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_readable = monroe_ionphoton_rtio_core_outputs_record3_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_seqn0 = monroe_ionphoton_rtio_core_outputs_record3_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record3_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address0 = monroe_ionphoton_rtio_core_outputs_record3_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data0 = monroe_ionphoton_rtio_core_outputs_record3_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record4_re = monroe_ionphoton_rtio_core_outputs_gates_record4_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_readable = monroe_ionphoton_rtio_core_outputs_record4_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_seqn0 = monroe_ionphoton_rtio_core_outputs_record4_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record4_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address0 = monroe_ionphoton_rtio_core_outputs_record4_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data0 = monroe_ionphoton_rtio_core_outputs_record4_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record5_re = monroe_ionphoton_rtio_core_outputs_gates_record5_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_readable = monroe_ionphoton_rtio_core_outputs_record5_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_seqn0 = monroe_ionphoton_rtio_core_outputs_record5_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record5_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address0 = monroe_ionphoton_rtio_core_outputs_record5_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data0 = monroe_ionphoton_rtio_core_outputs_record5_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record6_re = monroe_ionphoton_rtio_core_outputs_gates_record6_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_readable = monroe_ionphoton_rtio_core_outputs_record6_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_seqn0 = monroe_ionphoton_rtio_core_outputs_record6_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record6_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address0 = monroe_ionphoton_rtio_core_outputs_record6_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data0 = monroe_ionphoton_rtio_core_outputs_record6_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record7_re = monroe_ionphoton_rtio_core_outputs_gates_record7_re;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_readable = monroe_ionphoton_rtio_core_outputs_record7_readable;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_seqn0 = monroe_ionphoton_rtio_core_outputs_record7_seqn1;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel0 = monroe_ionphoton_rtio_core_outputs_record7_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_payload_timestamp = monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp1;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address0 = monroe_ionphoton_rtio_core_outputs_record7_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data0 = monroe_ionphoton_rtio_core_outputs_record7_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record0_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record0_valid;
assign monroe_ionphoton_rtio_core_outputs_record0_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record0_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record0_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record0_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record0_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record0_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record0_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record1_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record1_valid;
assign monroe_ionphoton_rtio_core_outputs_record1_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record1_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record1_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record1_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record1_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record1_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record1_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record2_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record2_valid;
assign monroe_ionphoton_rtio_core_outputs_record2_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record2_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record2_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record2_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record2_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record2_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record2_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record3_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record3_valid;
assign monroe_ionphoton_rtio_core_outputs_record3_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record3_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record3_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record3_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record3_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record3_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record3_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record4_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record4_valid;
assign monroe_ionphoton_rtio_core_outputs_record4_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record4_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record4_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record4_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record4_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record4_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record4_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record5_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record5_valid;
assign monroe_ionphoton_rtio_core_outputs_record5_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record5_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record5_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record5_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record5_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record5_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record5_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record6_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record6_valid;
assign monroe_ionphoton_rtio_core_outputs_record6_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record6_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record6_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record6_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record6_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record6_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record6_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data1;
assign monroe_ionphoton_rtio_core_outputs_record7_valid0 = monroe_ionphoton_rtio_core_outputs_gates_record7_valid;
assign monroe_ionphoton_rtio_core_outputs_record7_seqn2 = monroe_ionphoton_rtio_core_outputs_gates_record7_seqn1;
assign monroe_ionphoton_rtio_core_outputs_record7_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record7_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured = monroe_ionphoton_rtio_core_outputs_gates_record7_nondata_replace_occured;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_channel2 = monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel1;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0 = monroe_ionphoton_rtio_core_outputs_gates_record7_payload_fine_ts;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_address2 = monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address1;
assign monroe_ionphoton_rtio_core_outputs_record7_payload_data2 = monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data1;
assign monroe_ionphoton_rtio_core_cri_o_status = {monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_underflow, monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_wait};
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_seqn = monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_channel = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_address = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_data = monroe_ionphoton_rtio_core_cri_o_data;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp = monroe_ionphoton_rtio_core_cri_o_timestamp[63:3];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_plus_one = (monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane + 1'd1);
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_adr = monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation = monroe_ionphoton_rtio_core_outputs_lanedistributor_dat_r;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_min = ((monroe_ionphoton_rtio_core_outputs_lanedistributor_min_minus_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min = ((monroe_ionphoton_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min = ((monroe_ionphoton_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_last = ((monroe_ionphoton_rtio_core_outputs_lanedistributor_last_minus_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));

// synthesis translate_off
reg dummy_d_82;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen <= 3'd0;
	if ((monroe_ionphoton_rtio_core_outputs_lanedistributor_force_laneB | (~monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_last))) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen <= monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_plus_one;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_use_laneB <= 1'd1;
	end else begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen <= monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	end
// synthesis translate_off
	dummy_d_82 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_lane_min = (monroe_ionphoton_rtio_core_outputs_lanedistributor_use_laneB ? monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min : monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min);

// synthesis translate_off
reg dummy_d_83;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_do_underflow <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd0;
	if (((~monroe_ionphoton_rtio_core_outputs_lanedistributor_quash) & (monroe_ionphoton_rtio_core_cri_cmd == 1'd1))) begin
		if (monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_min) begin
			if (monroe_ionphoton_rtio_core_outputs_lanedistributor_timestamp_above_lane_min) begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write <= 1'd1;
			end else begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd1;
			end
		end else begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_do_underflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_83 <= dummy_s;
// synthesis translate_on
end
assign comb_lhs_array_muxed = monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write;

// synthesis translate_off
reg dummy_d_84;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_we <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_we <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen)
		1'd0: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_we <= comb_lhs_array_muxed;
		end
		1'd1: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_we <= comb_lhs_array_muxed;
		end
		2'd2: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_we <= comb_lhs_array_muxed;
		end
		2'd3: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_we <= comb_lhs_array_muxed;
		end
		3'd4: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_we <= comb_lhs_array_muxed;
		end
		3'd5: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_we <= comb_lhs_array_muxed;
		end
		3'd6: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_we <= comb_lhs_array_muxed;
		end
		default: begin
			monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_we <= comb_lhs_array_muxed;
		end
	endcase
// synthesis translate_off
	dummy_d_84 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp = ($signed({1'd0, monroe_ionphoton_rtio_core_cri_o_timestamp}) + (monroe_ionphoton_rtio_core_outputs_lanedistributor_compensation <<< 2'd3));

// synthesis translate_off
reg dummy_d_85;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_85 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_86;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_86 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_87;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_87 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_88;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_88 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_89;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_89 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_90;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_90 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_91;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_91 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_92;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= 64'd0;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_92 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable = comb_rhs_array_muxed8;
assign monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_wait = (~monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din = {{monroe_ionphoton_rtio_core_outputs_record0_payload_data0, monroe_ionphoton_rtio_core_outputs_record0_payload_address0, monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record0_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record0_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we = monroe_ionphoton_rtio_core_outputs_record0_we;
assign monroe_ionphoton_rtio_core_outputs_record0_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record0_payload_data1, monroe_ionphoton_rtio_core_outputs_record0_payload_address1, monroe_ionphoton_rtio_core_outputs_record0_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record0_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record0_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_dout;
assign monroe_ionphoton_rtio_core_outputs_record0_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_re = monroe_ionphoton_rtio_core_outputs_record0_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din = {{monroe_ionphoton_rtio_core_outputs_record1_payload_data0, monroe_ionphoton_rtio_core_outputs_record1_payload_address0, monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record1_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record1_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we = monroe_ionphoton_rtio_core_outputs_record1_we;
assign monroe_ionphoton_rtio_core_outputs_record1_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record1_payload_data1, monroe_ionphoton_rtio_core_outputs_record1_payload_address1, monroe_ionphoton_rtio_core_outputs_record1_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record1_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record1_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_dout;
assign monroe_ionphoton_rtio_core_outputs_record1_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_re = monroe_ionphoton_rtio_core_outputs_record1_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din = {{monroe_ionphoton_rtio_core_outputs_record2_payload_data0, monroe_ionphoton_rtio_core_outputs_record2_payload_address0, monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record2_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record2_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we = monroe_ionphoton_rtio_core_outputs_record2_we;
assign monroe_ionphoton_rtio_core_outputs_record2_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record2_payload_data1, monroe_ionphoton_rtio_core_outputs_record2_payload_address1, monroe_ionphoton_rtio_core_outputs_record2_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record2_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record2_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_dout;
assign monroe_ionphoton_rtio_core_outputs_record2_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_re = monroe_ionphoton_rtio_core_outputs_record2_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din = {{monroe_ionphoton_rtio_core_outputs_record3_payload_data0, monroe_ionphoton_rtio_core_outputs_record3_payload_address0, monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record3_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record3_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we = monroe_ionphoton_rtio_core_outputs_record3_we;
assign monroe_ionphoton_rtio_core_outputs_record3_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record3_payload_data1, monroe_ionphoton_rtio_core_outputs_record3_payload_address1, monroe_ionphoton_rtio_core_outputs_record3_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record3_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record3_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_dout;
assign monroe_ionphoton_rtio_core_outputs_record3_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_re = monroe_ionphoton_rtio_core_outputs_record3_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din = {{monroe_ionphoton_rtio_core_outputs_record4_payload_data0, monroe_ionphoton_rtio_core_outputs_record4_payload_address0, monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record4_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record4_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we = monroe_ionphoton_rtio_core_outputs_record4_we;
assign monroe_ionphoton_rtio_core_outputs_record4_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record4_payload_data1, monroe_ionphoton_rtio_core_outputs_record4_payload_address1, monroe_ionphoton_rtio_core_outputs_record4_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record4_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record4_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_dout;
assign monroe_ionphoton_rtio_core_outputs_record4_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_re = monroe_ionphoton_rtio_core_outputs_record4_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din = {{monroe_ionphoton_rtio_core_outputs_record5_payload_data0, monroe_ionphoton_rtio_core_outputs_record5_payload_address0, monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record5_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record5_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we = monroe_ionphoton_rtio_core_outputs_record5_we;
assign monroe_ionphoton_rtio_core_outputs_record5_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record5_payload_data1, monroe_ionphoton_rtio_core_outputs_record5_payload_address1, monroe_ionphoton_rtio_core_outputs_record5_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record5_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record5_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_dout;
assign monroe_ionphoton_rtio_core_outputs_record5_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_re = monroe_ionphoton_rtio_core_outputs_record5_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din = {{monroe_ionphoton_rtio_core_outputs_record6_payload_data0, monroe_ionphoton_rtio_core_outputs_record6_payload_address0, monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record6_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record6_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we = monroe_ionphoton_rtio_core_outputs_record6_we;
assign monroe_ionphoton_rtio_core_outputs_record6_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record6_payload_data1, monroe_ionphoton_rtio_core_outputs_record6_payload_address1, monroe_ionphoton_rtio_core_outputs_record6_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record6_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record6_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_dout;
assign monroe_ionphoton_rtio_core_outputs_record6_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_re = monroe_ionphoton_rtio_core_outputs_record6_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din = {{monroe_ionphoton_rtio_core_outputs_record7_payload_data0, monroe_ionphoton_rtio_core_outputs_record7_payload_address0, monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp0, monroe_ionphoton_rtio_core_outputs_record7_payload_channel0}, monroe_ionphoton_rtio_core_outputs_record7_seqn0};
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we = monroe_ionphoton_rtio_core_outputs_record7_we;
assign monroe_ionphoton_rtio_core_outputs_record7_writable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
assign {{monroe_ionphoton_rtio_core_outputs_record7_payload_data1, monroe_ionphoton_rtio_core_outputs_record7_payload_address1, monroe_ionphoton_rtio_core_outputs_record7_payload_timestamp1, monroe_ionphoton_rtio_core_outputs_record7_payload_channel1}, monroe_ionphoton_rtio_core_outputs_record7_seqn1} = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_dout;
assign monroe_ionphoton_rtio_core_outputs_record7_readable = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_re = monroe_ionphoton_rtio_core_outputs_record7_re;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_93;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_93 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_94;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_94 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_95;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_95 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_96;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_96 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_97;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_97 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_98;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_98 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_99;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_99 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_100;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_100 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_101;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_101 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_102;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_102 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_103;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_103 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_104;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_104 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_105;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_105 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_106;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_106 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable & monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable = (((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[7] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[7]) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[6] == monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[6])) | (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[5:0] != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[5:0]));
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q != monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_produce_rdomain);
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_we = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_adr = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[6:0];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout = monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;

// synthesis translate_off
reg dummy_d_107;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary;
	end
// synthesis translate_off
	dummy_d_107 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_108;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= 8'd0;
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary;
	end
// synthesis translate_off
	dummy_d_108 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next = (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary ^ monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[7:1]);
assign monroe_ionphoton_rtio_core_outputs_gates_record0_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record0_re = (monroe_ionphoton_rtio_core_outputs_gates_record0_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record1_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record1_re = (monroe_ionphoton_rtio_core_outputs_gates_record1_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record2_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record2_re = (monroe_ionphoton_rtio_core_outputs_gates_record2_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record3_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record3_re = (monroe_ionphoton_rtio_core_outputs_gates_record3_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record4_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record4_re = (monroe_ionphoton_rtio_core_outputs_gates_record4_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record5_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record5_re = (monroe_ionphoton_rtio_core_outputs_gates_record5_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record6_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record6_re = (monroe_ionphoton_rtio_core_outputs_gates_record6_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_gates_record7_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_nondata_replace_occured = 1'd0;
assign monroe_ionphoton_rtio_core_outputs_gates_record7_re = (monroe_ionphoton_rtio_core_outputs_gates_record7_payload_timestamp[63:3] == monroe_ionphoton_rtio_core_outputs_gates_coarse_timestamp);
assign monroe_ionphoton_rtio_core_outputs_memory0_adr = monroe_ionphoton_rtio_core_outputs_record40_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record0_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r0 & ((~monroe_ionphoton_rtio_core_outputs_memory0_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r0));
assign monroe_ionphoton_rtio_core_outputs_memory1_adr = monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record1_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r1 & ((~monroe_ionphoton_rtio_core_outputs_memory1_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r1));
assign monroe_ionphoton_rtio_core_outputs_memory2_adr = monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record2_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r2 & ((~monroe_ionphoton_rtio_core_outputs_memory2_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r2));
assign monroe_ionphoton_rtio_core_outputs_memory3_adr = monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record3_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r3 & ((~monroe_ionphoton_rtio_core_outputs_memory3_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r3));
assign monroe_ionphoton_rtio_core_outputs_memory4_adr = monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record4_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r4 & ((~monroe_ionphoton_rtio_core_outputs_memory4_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r4));
assign monroe_ionphoton_rtio_core_outputs_memory5_adr = monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record5_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r5 & ((~monroe_ionphoton_rtio_core_outputs_memory5_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r5));
assign monroe_ionphoton_rtio_core_outputs_memory6_adr = monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record6_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r6 & ((~monroe_ionphoton_rtio_core_outputs_memory6_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r6));
assign monroe_ionphoton_rtio_core_outputs_memory7_adr = monroe_ionphoton_rtio_core_outputs_record47_rec_payload_channel;
assign monroe_ionphoton_rtio_core_outputs_record7_collision = (monroe_ionphoton_rtio_core_outputs_replace_occured_r7 & ((~monroe_ionphoton_rtio_core_outputs_memory7_dat_r) | monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r7));
assign monroe_ionphoton_rtio_core_outputs_selected0 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected1 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected2 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected3 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected4 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected5 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected6 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected7 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 1'd0));
assign monroe_ionphoton_rtio_core_outputs_selected8 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected9 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected10 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected11 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected12 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected13 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected14 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected15 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 1'd1));
assign monroe_ionphoton_rtio_core_outputs_selected16 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected17 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected18 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected19 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected20 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected21 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected22 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected23 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 2'd2));
assign monroe_ionphoton_rtio_core_outputs_selected24 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected25 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected26 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected27 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected28 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected29 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected30 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected31 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 2'd3));
assign monroe_ionphoton_rtio_core_outputs_selected32 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected33 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected34 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected35 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected36 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected37 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected38 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected39 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 3'd4));
assign monroe_ionphoton_rtio_core_outputs_selected40 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected41 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected42 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected43 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected44 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected45 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected46 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected47 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 3'd5));
assign monroe_ionphoton_rtio_core_outputs_selected48 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected49 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected50 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected51 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected52 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected53 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected54 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected55 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 3'd6));
assign monroe_ionphoton_rtio_core_outputs_selected56 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected57 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected58 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected59 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected60 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected61 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected62 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected63 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 3'd7));
assign monroe_ionphoton_rtio_core_outputs_selected64 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected65 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected66 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected67 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected68 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected69 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected70 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected71 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd8));
assign monroe_ionphoton_rtio_core_outputs_selected72 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected73 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected74 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected75 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected76 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected77 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected78 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected79 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd9));
assign monroe_ionphoton_rtio_core_outputs_selected80 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected81 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected82 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected83 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected84 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected85 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected86 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected87 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd10));
assign monroe_ionphoton_rtio_core_outputs_selected88 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected89 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected90 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected91 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected92 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected93 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected94 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected95 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd11));
assign monroe_ionphoton_rtio_core_outputs_selected96 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected97 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected98 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected99 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected100 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected101 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected102 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected103 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd12));
assign monroe_ionphoton_rtio_core_outputs_selected104 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected105 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected106 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected107 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected108 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected109 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected110 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected111 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd13));
assign monroe_ionphoton_rtio_core_outputs_selected112 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected113 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected114 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected115 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected116 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected117 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected118 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected119 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd14));
assign monroe_ionphoton_rtio_core_outputs_selected120 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected121 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected122 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected123 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected124 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected125 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected126 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected127 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 4'd15));
assign monroe_ionphoton_rtio_core_outputs_selected128 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected129 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected130 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected131 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected132 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected133 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected134 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected135 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd16));
assign monroe_ionphoton_rtio_core_outputs_selected136 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected137 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected138 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected139 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected140 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected141 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected142 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected143 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd17));
assign monroe_ionphoton_rtio_core_outputs_selected144 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected145 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected146 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected147 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected148 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected149 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected150 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected151 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd18));
assign monroe_ionphoton_rtio_core_outputs_selected152 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected153 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected154 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected155 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected156 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected157 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected158 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected159 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd19));
assign monroe_ionphoton_rtio_core_outputs_selected160 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected161 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected162 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected163 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected164 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected165 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected166 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected167 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd20));
assign monroe_ionphoton_rtio_core_outputs_selected168 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected169 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected170 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected171 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected172 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected173 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected174 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected175 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd21));
assign monroe_ionphoton_rtio_core_outputs_selected176 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected177 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected178 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected179 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected180 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected181 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected182 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected183 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd22));
assign monroe_ionphoton_rtio_core_outputs_selected184 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected185 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected186 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected187 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected188 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected189 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected190 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected191 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd23));
assign monroe_ionphoton_rtio_core_outputs_selected192 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected193 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected194 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected195 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected196 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected197 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected198 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected199 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd24));
assign monroe_ionphoton_rtio_core_outputs_selected200 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected201 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected202 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected203 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected204 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected205 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected206 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected207 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd25));
assign monroe_ionphoton_rtio_core_outputs_selected208 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected209 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected210 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected211 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected212 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected213 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected214 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected215 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd26));
assign monroe_ionphoton_rtio_core_outputs_selected216 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected217 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected218 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected219 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected220 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected221 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected222 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected223 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd27));
assign monroe_ionphoton_rtio_core_outputs_selected224 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected225 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected226 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected227 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected228 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected229 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected230 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected231 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd28));
assign monroe_ionphoton_rtio_core_outputs_selected232 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected233 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected234 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected235 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected236 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected237 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected238 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected239 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd29));
assign monroe_ionphoton_rtio_core_outputs_selected240 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected241 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected242 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected243 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected244 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected245 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected246 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected247 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd30));
assign monroe_ionphoton_rtio_core_outputs_selected248 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected249 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected250 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected251 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected252 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected253 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected254 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected255 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 5'd31));
assign monroe_ionphoton_rtio_core_outputs_selected256 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected257 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected258 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected259 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected260 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected261 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected262 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected263 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 6'd32));
assign monroe_ionphoton_rtio_core_outputs_selected264 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected265 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected266 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected267 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected268 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected269 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected270 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected271 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 6'd33));
assign monroe_ionphoton_rtio_core_outputs_selected272 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected273 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected274 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected275 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected276 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected277 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected278 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected279 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 6'd34));
assign monroe_ionphoton_rtio_core_outputs_selected280 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected281 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected282 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected283 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected284 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected285 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected286 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected287 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 6'd35));
assign monroe_ionphoton_rtio_core_outputs_selected288 = ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision)) & (monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected289 = ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision)) & (monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected290 = ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision)) & (monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected291 = ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision)) & (monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected292 = ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision)) & (monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected293 = ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision)) & (monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected294 = ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision)) & (monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 == 6'd36));
assign monroe_ionphoton_rtio_core_outputs_selected295 = ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision)) & (monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 == 6'd36));

// synthesis translate_off
reg dummy_d_109;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference0 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record0_payload_channel2 != monroe_ionphoton_rtio_core_outputs_record1_payload_channel2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0 != monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record0_payload_address2 != monroe_ionphoton_rtio_core_outputs_record1_payload_address2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_109 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_110;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference1 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record2_payload_channel2 != monroe_ionphoton_rtio_core_outputs_record3_payload_channel2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0 != monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record2_payload_address2 != monroe_ionphoton_rtio_core_outputs_record3_payload_address2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_110 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_111;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference2 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record4_payload_channel2 != monroe_ionphoton_rtio_core_outputs_record5_payload_channel2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0 != monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record4_payload_address2 != monroe_ionphoton_rtio_core_outputs_record5_payload_address2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_111 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_112;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference3 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record6_payload_channel2 != monroe_ionphoton_rtio_core_outputs_record7_payload_channel2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0 != monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record6_payload_address2 != monroe_ionphoton_rtio_core_outputs_record7_payload_address2)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_112 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_113;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference4 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_113 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_114;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference5 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_114 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_115;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference6 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_115 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_116;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference7 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_116 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_117;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference8 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_117 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_118;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference9 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_118 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_119;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference10 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_119 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_120;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference11 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_120 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_121;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference12 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_121 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_122;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference13 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_122 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_123;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference14 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_123 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_124;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference15 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_124 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_125;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference16 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_125 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_126;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference17 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_126 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_127;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_outputs_nondata_difference18 <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel != monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts != monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address != monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address)) begin
		monroe_ionphoton_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_127 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_din = {monroe_ionphoton_rtio_core_inputs_record0_fifo_in_timestamp, monroe_ionphoton_rtio_core_inputs_record0_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record0_fifo_out_timestamp, monroe_ionphoton_rtio_core_inputs_record0_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
assign monroe_ionphoton_rtio_core_inputs_record0_fifo_in_data = inout_8x0_inout_8x0_iinterface0_data;
assign monroe_ionphoton_rtio_core_inputs_record0_fifo_in_timestamp = {monroe_ionphoton_rtio_tsc_coarse_ts, inout_8x0_inout_8x0_iinterface0_fine_ts};
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_we = inout_8x0_inout_8x0_iinterface0_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io0 = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_i = monroe_ionphoton_rtio_core_inputs_overflow_io0;
assign monroe_ionphoton_rtio_core_inputs_selected0 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 1'd0);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_re = ((monroe_ionphoton_rtio_core_inputs_selected0 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow0));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_din = {monroe_ionphoton_rtio_core_inputs_record1_fifo_in_timestamp, monroe_ionphoton_rtio_core_inputs_record1_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record1_fifo_out_timestamp, monroe_ionphoton_rtio_core_inputs_record1_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
assign monroe_ionphoton_rtio_core_inputs_record1_fifo_in_data = inout_8x1_inout_8x1_iinterface1_data;
assign monroe_ionphoton_rtio_core_inputs_record1_fifo_in_timestamp = {monroe_ionphoton_rtio_tsc_coarse_ts, inout_8x1_inout_8x1_iinterface1_fine_ts};
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_we = inout_8x1_inout_8x1_iinterface1_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io1 = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_i = monroe_ionphoton_rtio_core_inputs_overflow_io1;
assign monroe_ionphoton_rtio_core_inputs_selected1 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 1'd1);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_re = ((monroe_ionphoton_rtio_core_inputs_selected1 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow1));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_din = {monroe_ionphoton_rtio_core_inputs_record2_fifo_in_timestamp, monroe_ionphoton_rtio_core_inputs_record2_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record2_fifo_out_timestamp, monroe_ionphoton_rtio_core_inputs_record2_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
assign monroe_ionphoton_rtio_core_inputs_record2_fifo_in_data = inout_8x2_inout_8x2_iinterface2_data;
assign monroe_ionphoton_rtio_core_inputs_record2_fifo_in_timestamp = {monroe_ionphoton_rtio_tsc_coarse_ts, inout_8x2_inout_8x2_iinterface2_fine_ts};
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_we = inout_8x2_inout_8x2_iinterface2_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io2 = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_i = monroe_ionphoton_rtio_core_inputs_overflow_io2;
assign monroe_ionphoton_rtio_core_inputs_selected2 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 2'd2);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_re = ((monroe_ionphoton_rtio_core_inputs_selected2 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow2));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_din = {monroe_ionphoton_rtio_core_inputs_record3_fifo_in_timestamp, monroe_ionphoton_rtio_core_inputs_record3_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record3_fifo_out_timestamp, monroe_ionphoton_rtio_core_inputs_record3_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
assign monroe_ionphoton_rtio_core_inputs_record3_fifo_in_data = inout_8x3_inout_8x3_iinterface3_data;
assign monroe_ionphoton_rtio_core_inputs_record3_fifo_in_timestamp = {monroe_ionphoton_rtio_tsc_coarse_ts, inout_8x3_inout_8x3_iinterface3_fine_ts};
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_we = inout_8x3_inout_8x3_iinterface3_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io3 = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_i = monroe_ionphoton_rtio_core_inputs_overflow_io3;
assign monroe_ionphoton_rtio_core_inputs_selected3 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 2'd3);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_re = ((monroe_ionphoton_rtio_core_inputs_selected3 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow3));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_din = {monroe_ionphoton_rtio_core_inputs_record4_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record4_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
assign monroe_ionphoton_rtio_core_inputs_record4_fifo_in_data = spimaster0_iinterface0_data;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_we = spimaster0_iinterface0_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io4 = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_i = monroe_ionphoton_rtio_core_inputs_overflow_io4;
assign monroe_ionphoton_rtio_core_inputs_selected4 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 5'd16);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_re = ((monroe_ionphoton_rtio_core_inputs_selected4 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow4));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_din = {monroe_ionphoton_rtio_core_inputs_record5_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record5_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
assign monroe_ionphoton_rtio_core_inputs_record5_fifo_in_data = spimaster1_iinterface1_data;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_we = spimaster1_iinterface1_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io5 = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_i = monroe_ionphoton_rtio_core_inputs_overflow_io5;
assign monroe_ionphoton_rtio_core_inputs_selected5 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 5'd22);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_re = ((monroe_ionphoton_rtio_core_inputs_selected5 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow5));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_din = {monroe_ionphoton_rtio_core_inputs_record6_fifo_in_data};
assign {monroe_ionphoton_rtio_core_inputs_record6_fifo_out_data} = monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
assign monroe_ionphoton_rtio_core_inputs_record6_fifo_in_data = spimaster2_iinterface2_data;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_we = spimaster2_iinterface2_stb;
assign monroe_ionphoton_rtio_core_inputs_overflow_io6 = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_we & (~monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_writable));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_i = monroe_ionphoton_rtio_core_inputs_overflow_io6;
assign monroe_ionphoton_rtio_core_inputs_selected6 = (monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 5'd28);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_re = ((monroe_ionphoton_rtio_core_inputs_selected6 & monroe_ionphoton_rtio_core_inputs_i_ack) & (~monroe_ionphoton_rtio_core_inputs_overflow6));
assign monroe_ionphoton_rtio_core_inputs_i_status_raw = comb_rhs_array_muxed9;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q[6] == monroe_ionphoton_rtio_core_inputs_asyncfifo0_consume_wdomain[6]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q[5] == monroe_ionphoton_rtio_core_inputs_asyncfifo0_consume_wdomain[5])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q[4:0] != monroe_ionphoton_rtio_core_inputs_asyncfifo0_consume_wdomain[4:0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q != monroe_ionphoton_rtio_core_inputs_asyncfifo0_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_128;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_128 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_129;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_129 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[6:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer0_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer0_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_o = monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q[6] == monroe_ionphoton_rtio_core_inputs_asyncfifo1_consume_wdomain[6]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q[5] == monroe_ionphoton_rtio_core_inputs_asyncfifo1_consume_wdomain[5])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q[4:0] != monroe_ionphoton_rtio_core_inputs_asyncfifo1_consume_wdomain[4:0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q != monroe_ionphoton_rtio_core_inputs_asyncfifo1_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_130;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_130 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_131;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_131 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[6:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer1_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer1_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_o = monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q[6] == monroe_ionphoton_rtio_core_inputs_asyncfifo2_consume_wdomain[6]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q[5] == monroe_ionphoton_rtio_core_inputs_asyncfifo2_consume_wdomain[5])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q[4:0] != monroe_ionphoton_rtio_core_inputs_asyncfifo2_consume_wdomain[4:0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q != monroe_ionphoton_rtio_core_inputs_asyncfifo2_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_132;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_132 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_133;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_133 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[6:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer2_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer2_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_o = monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q[6] == monroe_ionphoton_rtio_core_inputs_asyncfifo3_consume_wdomain[6]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q[5] == monroe_ionphoton_rtio_core_inputs_asyncfifo3_consume_wdomain[5])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q[4:0] != monroe_ionphoton_rtio_core_inputs_asyncfifo3_consume_wdomain[4:0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q != monroe_ionphoton_rtio_core_inputs_asyncfifo3_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[5:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_134;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_134 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_135;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= 7'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_135 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[6:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer3_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer3_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_o = monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q[2] == monroe_ionphoton_rtio_core_inputs_asyncfifo4_consume_wdomain[2]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q[1] == monroe_ionphoton_rtio_core_inputs_asyncfifo4_consume_wdomain[1])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q[0] != monroe_ionphoton_rtio_core_inputs_asyncfifo4_consume_wdomain[0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q != monroe_ionphoton_rtio_core_inputs_asyncfifo4_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_136;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_136 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_137;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_137 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[2:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer4_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer4_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_o = monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q[2] == monroe_ionphoton_rtio_core_inputs_asyncfifo5_consume_wdomain[2]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q[1] == monroe_ionphoton_rtio_core_inputs_asyncfifo5_consume_wdomain[1])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q[0] != monroe_ionphoton_rtio_core_inputs_asyncfifo5_consume_wdomain[0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q != monroe_ionphoton_rtio_core_inputs_asyncfifo5_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_138;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_138 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_139;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_139 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[2:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer5_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer5_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_o = monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_writable & monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_we);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_ce = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_re);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_writable = (((monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q[2] == monroe_ionphoton_rtio_core_inputs_asyncfifo6_consume_wdomain[2]) | (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q[1] == monroe_ionphoton_rtio_core_inputs_asyncfifo6_consume_wdomain[1])) | (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q[0] != monroe_ionphoton_rtio_core_inputs_asyncfifo6_consume_wdomain[0]));
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_readable = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q != monroe_ionphoton_rtio_core_inputs_asyncfifo6_produce_rdomain);
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_dat_w = monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_we = monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_ce;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_adr = monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[1:0];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_dout = monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_140;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_140 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_141;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= 3'd0;
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_ce) begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_binary + 1'd1);
	end else begin
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_141 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next = (monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary ^ monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[2:1]);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_i = (monroe_ionphoton_rtio_core_inputs_blindtransfer6_i & (~monroe_ionphoton_rtio_core_inputs_blindtransfer6_blind));
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_i = monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_o = monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_o;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_o = (monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_i = (monroe_ionphoton_rtio_core_o_collision_sync_i & (~monroe_ionphoton_rtio_core_o_collision_sync_blind));
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_i = monroe_ionphoton_rtio_core_o_collision_sync_ps_o;
assign monroe_ionphoton_rtio_core_o_collision_sync_o = monroe_ionphoton_rtio_core_o_collision_sync_ps_o;
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_o = (monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o ^ monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_o = (monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_i = (monroe_ionphoton_rtio_core_o_busy_sync_i & (~monroe_ionphoton_rtio_core_o_busy_sync_blind));
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_i = monroe_ionphoton_rtio_core_o_busy_sync_ps_o;
assign monroe_ionphoton_rtio_core_o_busy_sync_o = monroe_ionphoton_rtio_core_o_busy_sync_ps_o;
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_o = (monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o ^ monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o_r);
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_o = (monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o ^ monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o_r);
assign monroe_ionphoton_rtio_now_hi_w = monroe_ionphoton_rtio_now[63:32];
assign monroe_ionphoton_rtio_now_lo_w = monroe_ionphoton_rtio_now[31:0];

// synthesis translate_off
reg dummy_d_142;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_cri_cmd <= 2'd0;
	monroe_ionphoton_rtio_cri_cmd <= 1'd0;
	if (monroe_ionphoton_rtio_o_data_re) begin
		monroe_ionphoton_rtio_cri_cmd <= 1'd1;
	end
	if (monroe_ionphoton_rtio_i_timeout_re) begin
		monroe_ionphoton_rtio_cri_cmd <= 2'd2;
	end
// synthesis translate_off
	dummy_d_142 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_cri_chan_sel = monroe_ionphoton_rtio_target_storage[31:8];
assign monroe_ionphoton_rtio_cri_o_timestamp = monroe_ionphoton_rtio_now;
assign monroe_ionphoton_rtio_cri_o_data = monroe_ionphoton_rtio_o_data_storage;
assign monroe_ionphoton_rtio_cri_o_address = monroe_ionphoton_rtio_target_storage[7:0];
assign monroe_ionphoton_rtio_o_status_status = monroe_ionphoton_rtio_cri_o_status;
assign monroe_ionphoton_rtio_cri_i_timeout = monroe_ionphoton_rtio_i_timeout_storage;
assign monroe_ionphoton_rtio_i_data_status = monroe_ionphoton_rtio_cri_i_data;
assign monroe_ionphoton_rtio_i_timestamp_status = monroe_ionphoton_rtio_cri_i_timestamp;
assign monroe_ionphoton_rtio_i_status_status = monroe_ionphoton_rtio_cri_i_status;
assign monroe_ionphoton_rtio_o_data_dat_w = 1'd0;
assign monroe_ionphoton_rtio_o_data_we = monroe_ionphoton_rtio_target_re;
assign monroe_ionphoton_dma_rawslicer_sink_stb = monroe_ionphoton_dma_dma_source_stb;
assign monroe_ionphoton_dma_dma_source_ack = monroe_ionphoton_dma_rawslicer_sink_ack;
assign monroe_ionphoton_dma_rawslicer_sink_eop = monroe_ionphoton_dma_dma_source_eop;
assign monroe_ionphoton_dma_rawslicer_sink_payload_data = monroe_ionphoton_dma_dma_source_payload_data;
assign monroe_ionphoton_dma_time_offset_sink_stb = monroe_ionphoton_dma_record_converter_source_stb;
assign monroe_ionphoton_dma_record_converter_source_ack = monroe_ionphoton_dma_time_offset_sink_ack;
assign monroe_ionphoton_dma_time_offset_sink_eop = monroe_ionphoton_dma_record_converter_source_eop;
assign monroe_ionphoton_dma_time_offset_sink_payload_length = monroe_ionphoton_dma_record_converter_source_payload_length;
assign monroe_ionphoton_dma_time_offset_sink_payload_channel = monroe_ionphoton_dma_record_converter_source_payload_channel;
assign monroe_ionphoton_dma_time_offset_sink_payload_timestamp = monroe_ionphoton_dma_record_converter_source_payload_timestamp;
assign monroe_ionphoton_dma_time_offset_sink_payload_address = monroe_ionphoton_dma_record_converter_source_payload_address;
assign monroe_ionphoton_dma_time_offset_sink_payload_data = monroe_ionphoton_dma_record_converter_source_payload_data;
assign monroe_ionphoton_dma_cri_master_sink_stb = monroe_ionphoton_dma_time_offset_source_stb;
assign monroe_ionphoton_dma_time_offset_source_ack = monroe_ionphoton_dma_cri_master_sink_ack;
assign monroe_ionphoton_dma_cri_master_sink_eop = monroe_ionphoton_dma_time_offset_source_eop;
assign monroe_ionphoton_dma_cri_master_sink_payload_length = monroe_ionphoton_dma_time_offset_source_payload_length;
assign monroe_ionphoton_dma_cri_master_sink_payload_channel = monroe_ionphoton_dma_time_offset_source_payload_channel;
assign monroe_ionphoton_dma_cri_master_sink_payload_timestamp = monroe_ionphoton_dma_time_offset_source_payload_timestamp;
assign monroe_ionphoton_dma_cri_master_sink_payload_address = monroe_ionphoton_dma_time_offset_source_payload_address;
assign monroe_ionphoton_dma_cri_master_sink_payload_data = monroe_ionphoton_dma_time_offset_source_payload_data;
assign monroe_ionphoton_dma_dma_bus_stb = (monroe_ionphoton_dma_dma_sink_stb & ((~monroe_ionphoton_dma_dma_data_reg_loaded) | monroe_ionphoton_dma_dma_source_ack));
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_cyc = monroe_ionphoton_dma_dma_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_stb = monroe_ionphoton_dma_dma_bus_stb;
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_adr = monroe_ionphoton_dma_dma_sink_payload_address;
assign monroe_ionphoton_dma_dma_sink_ack = monroe_ionphoton_monroe_ionphoton_interface0_bus_ack;
assign monroe_ionphoton_dma_dma_source_stb = monroe_ionphoton_dma_dma_data_reg_loaded;
assign monroe_ionphoton_dma_rawslicer_source = monroe_ionphoton_dma_rawslicer_buf[615:0];

// synthesis translate_off
reg dummy_d_143;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_dma_rawslicer_sink_ack <= 1'd0;
	monroe_ionphoton_dma_rawslicer_source_stb <= 1'd0;
	monroe_ionphoton_dma_rawslicer_flush_done <= 1'd0;
	monroe_ionphoton_dma_rawslicer_next_level <= 7'd0;
	monroe_ionphoton_dma_rawslicer_load_buf <= 1'd0;
	monroe_ionphoton_dma_rawslicer_shift_buf <= 1'd0;
	clockdomainsrenamer_resetinserter_next_state <= 2'd0;
	monroe_ionphoton_dma_rawslicer_next_level <= monroe_ionphoton_dma_rawslicer_level;
	clockdomainsrenamer_resetinserter_next_state <= clockdomainsrenamer_resetinserter_state;
	case (clockdomainsrenamer_resetinserter_state)
		1'd1: begin
			monroe_ionphoton_dma_rawslicer_source_stb <= 1'd1;
			monroe_ionphoton_dma_rawslicer_shift_buf <= 1'd1;
			monroe_ionphoton_dma_rawslicer_next_level <= (monroe_ionphoton_dma_rawslicer_level - monroe_ionphoton_dma_rawslicer_source_consume);
			if ((monroe_ionphoton_dma_rawslicer_next_level < 7'd77)) begin
				clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
			if (monroe_ionphoton_dma_rawslicer_flush) begin
				clockdomainsrenamer_resetinserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			monroe_ionphoton_dma_rawslicer_next_level <= 1'd0;
			monroe_ionphoton_dma_rawslicer_sink_ack <= 1'd1;
			if ((monroe_ionphoton_dma_rawslicer_sink_stb & monroe_ionphoton_dma_rawslicer_sink_eop)) begin
				monroe_ionphoton_dma_rawslicer_flush_done <= 1'd1;
				clockdomainsrenamer_resetinserter_next_state <= 1'd0;
			end
		end
		default: begin
			monroe_ionphoton_dma_rawslicer_sink_ack <= 1'd1;
			monroe_ionphoton_dma_rawslicer_load_buf <= 1'd1;
			if (monroe_ionphoton_dma_rawslicer_sink_stb) begin
				monroe_ionphoton_dma_rawslicer_next_level <= (monroe_ionphoton_dma_rawslicer_level + 5'd16);
			end
			if ((monroe_ionphoton_dma_rawslicer_next_level >= 7'd77)) begin
				clockdomainsrenamer_resetinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_143 <= dummy_s;
// synthesis translate_on
end
assign {monroe_ionphoton_dma_record_converter_record_raw_data, monroe_ionphoton_dma_record_converter_record_raw_address, monroe_ionphoton_dma_record_converter_record_raw_timestamp, monroe_ionphoton_dma_record_converter_record_raw_channel, monroe_ionphoton_dma_record_converter_record_raw_length} = monroe_ionphoton_dma_rawslicer_source;
assign monroe_ionphoton_dma_record_converter_source_payload_channel = monroe_ionphoton_dma_record_converter_record_raw_channel;
assign monroe_ionphoton_dma_record_converter_source_payload_timestamp = monroe_ionphoton_dma_record_converter_record_raw_timestamp;
assign monroe_ionphoton_dma_record_converter_source_payload_address = monroe_ionphoton_dma_record_converter_record_raw_address;

// synthesis translate_off
reg dummy_d_144;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_dma_record_converter_source_payload_data <= 512'd0;
	case (monroe_ionphoton_dma_record_converter_record_raw_length)
		4'd14: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[7:0];
		end
		4'd15: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[15:0];
		end
		5'd16: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[23:0];
		end
		5'd17: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[31:0];
		end
		5'd18: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[39:0];
		end
		5'd19: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[47:0];
		end
		5'd20: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[55:0];
		end
		5'd21: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[63:0];
		end
		5'd22: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[71:0];
		end
		5'd23: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[79:0];
		end
		5'd24: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[87:0];
		end
		5'd25: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[95:0];
		end
		5'd26: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[103:0];
		end
		5'd27: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[111:0];
		end
		5'd28: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[119:0];
		end
		5'd29: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[127:0];
		end
		5'd30: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[135:0];
		end
		5'd31: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[143:0];
		end
		6'd32: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[151:0];
		end
		6'd33: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[159:0];
		end
		6'd34: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[167:0];
		end
		6'd35: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[175:0];
		end
		6'd36: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[183:0];
		end
		6'd37: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[191:0];
		end
		6'd38: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[199:0];
		end
		6'd39: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[207:0];
		end
		6'd40: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[215:0];
		end
		6'd41: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[223:0];
		end
		6'd42: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[231:0];
		end
		6'd43: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[239:0];
		end
		6'd44: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[247:0];
		end
		6'd45: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[255:0];
		end
		6'd46: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[263:0];
		end
		6'd47: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[271:0];
		end
		6'd48: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[279:0];
		end
		6'd49: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[287:0];
		end
		6'd50: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[295:0];
		end
		6'd51: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[303:0];
		end
		6'd52: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[311:0];
		end
		6'd53: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[319:0];
		end
		6'd54: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[327:0];
		end
		6'd55: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[335:0];
		end
		6'd56: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[343:0];
		end
		6'd57: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[351:0];
		end
		6'd58: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[359:0];
		end
		6'd59: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[367:0];
		end
		6'd60: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[375:0];
		end
		6'd61: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[383:0];
		end
		6'd62: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[391:0];
		end
		6'd63: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[399:0];
		end
		7'd64: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[407:0];
		end
		7'd65: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[415:0];
		end
		7'd66: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[423:0];
		end
		7'd67: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[431:0];
		end
		7'd68: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[439:0];
		end
		7'd69: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[447:0];
		end
		7'd70: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[455:0];
		end
		7'd71: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[463:0];
		end
		7'd72: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[471:0];
		end
		7'd73: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[479:0];
		end
		7'd74: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[487:0];
		end
		7'd75: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[495:0];
		end
		7'd76: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[503:0];
		end
		7'd77: begin
			monroe_ionphoton_dma_record_converter_source_payload_data <= monroe_ionphoton_dma_record_converter_record_raw_data[511:0];
		end
	endcase
// synthesis translate_off
	dummy_d_144 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_145;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_dma_rawslicer_source_consume <= 7'd0;
	monroe_ionphoton_dma_rawslicer_flush <= 1'd0;
	monroe_ionphoton_dma_record_converter_source_stb <= 1'd0;
	monroe_ionphoton_dma_record_converter_source_eop <= 1'd0;
	monroe_ionphoton_dma_record_converter_end_marker_found <= 1'd0;
	clockdomainsrenamer_recordconverter_next_state <= 2'd0;
	clockdomainsrenamer_recordconverter_next_state <= clockdomainsrenamer_recordconverter_state;
	case (clockdomainsrenamer_recordconverter_state)
		1'd1: begin
			monroe_ionphoton_dma_record_converter_end_marker_found <= 1'd1;
			if (monroe_ionphoton_dma_record_converter_flush) begin
				monroe_ionphoton_dma_rawslicer_flush <= 1'd1;
				clockdomainsrenamer_recordconverter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (monroe_ionphoton_dma_rawslicer_flush_done) begin
				clockdomainsrenamer_recordconverter_next_state <= 2'd3;
			end
		end
		2'd3: begin
			monroe_ionphoton_dma_record_converter_source_eop <= 1'd1;
			monroe_ionphoton_dma_record_converter_source_stb <= 1'd1;
			if (monroe_ionphoton_dma_record_converter_source_ack) begin
				clockdomainsrenamer_recordconverter_next_state <= 1'd0;
			end
		end
		default: begin
			if (monroe_ionphoton_dma_rawslicer_source_stb) begin
				if ((monroe_ionphoton_dma_record_converter_record_raw_length == 1'd0)) begin
					clockdomainsrenamer_recordconverter_next_state <= 1'd1;
				end else begin
					monroe_ionphoton_dma_record_converter_source_stb <= 1'd1;
				end
			end
			if (monroe_ionphoton_dma_record_converter_source_ack) begin
				monroe_ionphoton_dma_rawslicer_source_consume <= monroe_ionphoton_dma_record_converter_record_raw_length;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_145 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_dma_time_offset_sink_ack = (~monroe_ionphoton_dma_time_offset_source_stb);
assign monroe_ionphoton_dma_cri_master_cri_chan_sel = monroe_ionphoton_dma_cri_master_sink_payload_channel;
assign monroe_ionphoton_dma_cri_master_cri_o_timestamp = monroe_ionphoton_dma_cri_master_sink_payload_timestamp;
assign monroe_ionphoton_dma_cri_master_cri_o_address = monroe_ionphoton_dma_cri_master_sink_payload_address;
assign monroe_ionphoton_dma_cri_master_cri_o_data = monroe_ionphoton_dma_cri_master_sink_payload_data;

// synthesis translate_off
reg dummy_d_146;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_dma_cri_master_sink_ack <= 1'd0;
	monroe_ionphoton_dma_cri_master_cri_cmd <= 2'd0;
	monroe_ionphoton_dma_cri_master_busy <= 1'd0;
	monroe_ionphoton_dma_cri_master_underflow_trigger <= 1'd0;
	monroe_ionphoton_dma_cri_master_link_error_trigger <= 1'd0;
	clockdomainsrenamer_crimaster_next_state <= 3'd0;
	clockdomainsrenamer_crimaster_next_state <= clockdomainsrenamer_crimaster_state;
	case (clockdomainsrenamer_crimaster_state)
		1'd1: begin
			monroe_ionphoton_dma_cri_master_busy <= 1'd1;
			monroe_ionphoton_dma_cri_master_cri_cmd <= 1'd1;
			clockdomainsrenamer_crimaster_next_state <= 2'd2;
		end
		2'd2: begin
			monroe_ionphoton_dma_cri_master_busy <= 1'd1;
			if ((monroe_ionphoton_dma_cri_master_cri_o_status == 1'd0)) begin
				monroe_ionphoton_dma_cri_master_sink_ack <= 1'd1;
				clockdomainsrenamer_crimaster_next_state <= 1'd0;
			end
			if (monroe_ionphoton_dma_cri_master_cri_o_status[1]) begin
				clockdomainsrenamer_crimaster_next_state <= 2'd3;
			end
			if (monroe_ionphoton_dma_cri_master_cri_o_status[2]) begin
				clockdomainsrenamer_crimaster_next_state <= 3'd4;
			end
		end
		2'd3: begin
			monroe_ionphoton_dma_cri_master_busy <= 1'd1;
			monroe_ionphoton_dma_cri_master_underflow_trigger <= 1'd1;
			monroe_ionphoton_dma_cri_master_sink_ack <= 1'd1;
			clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		3'd4: begin
			monroe_ionphoton_dma_cri_master_busy <= 1'd1;
			monroe_ionphoton_dma_cri_master_link_error_trigger <= 1'd1;
			monroe_ionphoton_dma_cri_master_sink_ack <= 1'd1;
			clockdomainsrenamer_crimaster_next_state <= 1'd0;
		end
		default: begin
			if ((monroe_ionphoton_dma_cri_master_error_w == 1'd0)) begin
				if (monroe_ionphoton_dma_cri_master_sink_stb) begin
					if (monroe_ionphoton_dma_cri_master_sink_eop) begin
						monroe_ionphoton_dma_cri_master_sink_ack <= 1'd1;
					end else begin
						clockdomainsrenamer_crimaster_next_state <= 1'd1;
					end
				end
			end else begin
				monroe_ionphoton_dma_cri_master_sink_ack <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_146 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_147;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_dma_enable_enable_w <= 1'd0;
	monroe_ionphoton_dma_flow_enable <= 1'd0;
	monroe_ionphoton_dma_record_converter_flush <= 1'd0;
	clockdomainsrenamer_fsm_next_state <= 3'd0;
	clockdomainsrenamer_fsm_next_state <= clockdomainsrenamer_fsm_state;
	case (clockdomainsrenamer_fsm_state)
		1'd1: begin
			monroe_ionphoton_dma_enable_enable_w <= 1'd1;
			monroe_ionphoton_dma_flow_enable <= 1'd1;
			if (monroe_ionphoton_dma_record_converter_end_marker_found) begin
				clockdomainsrenamer_fsm_next_state <= 2'd2;
			end
		end
		2'd2: begin
			monroe_ionphoton_dma_enable_enable_w <= 1'd1;
			monroe_ionphoton_dma_record_converter_flush <= 1'd1;
			clockdomainsrenamer_fsm_next_state <= 2'd3;
		end
		2'd3: begin
			monroe_ionphoton_dma_enable_enable_w <= 1'd1;
			if (((monroe_ionphoton_dma_cri_master_sink_stb & monroe_ionphoton_dma_cri_master_sink_ack) & monroe_ionphoton_dma_cri_master_sink_eop)) begin
				clockdomainsrenamer_fsm_next_state <= 3'd4;
			end
		end
		3'd4: begin
			monroe_ionphoton_dma_enable_enable_w <= 1'd1;
			if ((~monroe_ionphoton_dma_cri_master_busy)) begin
				clockdomainsrenamer_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			if (monroe_ionphoton_dma_enable_enable_re) begin
				clockdomainsrenamer_fsm_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_147 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_csrbank0_target0_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_target0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 1'd0));
assign monroe_ionphoton_rtio_now_hi_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_rtio_now_hi_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 1'd1));
assign monroe_ionphoton_rtio_now_lo_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_rtio_now_lo_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 2'd3));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 3'd4));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 3'd5));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 3'd6));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 3'd7));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd8));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd9));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd10));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd11));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd12));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd13));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd14));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 4'd15));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd16));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd17));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd18));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[2:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd19));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd20));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd21));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd22));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd23));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd24));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[3:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd25));
assign monroe_ionphoton_rtio_i_overflow_reset_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[0];
assign monroe_ionphoton_rtio_i_overflow_reset_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd26));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd27));
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd28));
assign monroe_ionphoton_rtio_counter_update_r = monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_w[0];
assign monroe_ionphoton_rtio_counter_update_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0] == 5'd29));
assign monroe_ionphoton_rtio_target_storage = monroe_ionphoton_rtio_target_storage_full[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_target0_w = monroe_ionphoton_rtio_target_storage_full[31:0];
assign monroe_ionphoton_rtio_o_data_storage = monroe_ionphoton_rtio_o_data_storage_full[511:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_w = monroe_ionphoton_rtio_o_data_storage_full[511:480];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_w = monroe_ionphoton_rtio_o_data_storage_full[479:448];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_w = monroe_ionphoton_rtio_o_data_storage_full[447:416];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_w = monroe_ionphoton_rtio_o_data_storage_full[415:384];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_w = monroe_ionphoton_rtio_o_data_storage_full[383:352];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_w = monroe_ionphoton_rtio_o_data_storage_full[351:320];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_w = monroe_ionphoton_rtio_o_data_storage_full[319:288];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_w = monroe_ionphoton_rtio_o_data_storage_full[287:256];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_w = monroe_ionphoton_rtio_o_data_storage_full[255:224];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_w = monroe_ionphoton_rtio_o_data_storage_full[223:192];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_w = monroe_ionphoton_rtio_o_data_storage_full[191:160];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_w = monroe_ionphoton_rtio_o_data_storage_full[159:128];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_w = monroe_ionphoton_rtio_o_data_storage_full[127:96];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_w = monroe_ionphoton_rtio_o_data_storage_full[95:64];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_w = monroe_ionphoton_rtio_o_data_storage_full[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_w = monroe_ionphoton_rtio_o_data_storage_full[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_w = monroe_ionphoton_rtio_o_status_status[2:0];
assign monroe_ionphoton_rtio_i_timeout_storage = monroe_ionphoton_rtio_i_timeout_storage_full[63:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_w = monroe_ionphoton_rtio_i_timeout_storage_full[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_w = monroe_ionphoton_rtio_i_timeout_storage_full[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_w = monroe_ionphoton_rtio_i_data_status[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_w = monroe_ionphoton_rtio_i_timestamp_status[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_w = monroe_ionphoton_rtio_i_timestamp_status[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_w = monroe_ionphoton_rtio_i_status_status[3:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_w = monroe_ionphoton_rtio_counter_status[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_w = monroe_ionphoton_rtio_counter_status[31:0];
assign monroe_ionphoton_dma_enable_enable_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[0];
assign monroe_ionphoton_dma_enable_enable_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[1:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 2'd3));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 3'd4));
assign monroe_ionphoton_dma_cri_master_error_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[1:0];
assign monroe_ionphoton_dma_cri_master_error_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 3'd5));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[23:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 3'd6));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 3'd7));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 4'd8));
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_r = monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_w[15:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0] == 4'd9));
assign monroe_ionphoton_dma_dma_storage = monroe_ionphoton_dma_dma_storage_full[33:4];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_w = monroe_ionphoton_dma_dma_storage_full[33:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_w = {monroe_ionphoton_dma_dma_storage_full[31:4], {28{1'd0}}};
assign monroe_ionphoton_dma_time_offset_storage = monroe_ionphoton_dma_time_offset_storage_full[63:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_w = monroe_ionphoton_dma_time_offset_storage_full[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_w = monroe_ionphoton_dma_time_offset_storage_full[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_w = monroe_ionphoton_dma_cri_master_error_channel_status[23:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_w = monroe_ionphoton_dma_cri_master_error_timestamp_status[63:32];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_w = monroe_ionphoton_dma_cri_master_error_timestamp_status[31:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_w = monroe_ionphoton_dma_cri_master_error_address_status[15:0];
assign monroe_ionphoton_cri_con_shared_cmd = comb_rhs_array_muxed10;
assign monroe_ionphoton_cri_con_shared_chan_sel = comb_rhs_array_muxed11;
assign monroe_ionphoton_cri_con_shared_o_timestamp = comb_rhs_array_muxed12;
assign monroe_ionphoton_cri_con_shared_o_data = comb_rhs_array_muxed13;
assign monroe_ionphoton_cri_con_shared_o_address = comb_rhs_array_muxed14;
assign monroe_ionphoton_cri_con_shared_i_timeout = comb_rhs_array_muxed15;
assign monroe_ionphoton_rtio_cri_o_status = monroe_ionphoton_cri_con_shared_o_status;
assign monroe_ionphoton_dma_cri_master_cri_o_status = monroe_ionphoton_cri_con_shared_o_status;
assign monroe_ionphoton_rtio_cri_o_buffer_space_valid = monroe_ionphoton_cri_con_shared_o_buffer_space_valid;
assign monroe_ionphoton_dma_cri_master_cri_o_buffer_space_valid = monroe_ionphoton_cri_con_shared_o_buffer_space_valid;
assign monroe_ionphoton_rtio_cri_o_buffer_space = monroe_ionphoton_cri_con_shared_o_buffer_space;
assign monroe_ionphoton_dma_cri_master_cri_o_buffer_space = monroe_ionphoton_cri_con_shared_o_buffer_space;
assign monroe_ionphoton_rtio_cri_i_data = monroe_ionphoton_cri_con_shared_i_data;
assign monroe_ionphoton_dma_cri_master_cri_i_data = monroe_ionphoton_cri_con_shared_i_data;
assign monroe_ionphoton_rtio_cri_i_timestamp = monroe_ionphoton_cri_con_shared_i_timestamp;
assign monroe_ionphoton_dma_cri_master_cri_i_timestamp = monroe_ionphoton_cri_con_shared_i_timestamp;
assign monroe_ionphoton_rtio_cri_i_status = monroe_ionphoton_cri_con_shared_i_status;
assign monroe_ionphoton_dma_cri_master_cri_i_status = monroe_ionphoton_cri_con_shared_i_status;
assign monroe_ionphoton_rtio_core_cri_chan_sel = monroe_ionphoton_cri_con_shared_chan_sel;
assign monroe_ionphoton_rtio_core_cri_o_timestamp = monroe_ionphoton_cri_con_shared_o_timestamp;
assign monroe_ionphoton_rtio_core_cri_o_data = monroe_ionphoton_cri_con_shared_o_data;
assign monroe_ionphoton_rtio_core_cri_o_address = monroe_ionphoton_cri_con_shared_o_address;
assign monroe_ionphoton_rtio_core_cri_i_timeout = monroe_ionphoton_cri_con_shared_i_timeout;

// synthesis translate_off
reg dummy_d_148;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_core_cri_cmd <= 2'd0;
	if ((monroe_ionphoton_cri_con_selected == 1'd0)) begin
		monroe_ionphoton_rtio_core_cri_cmd <= monroe_ionphoton_cri_con_shared_cmd;
	end
// synthesis translate_off
	dummy_d_148 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_149;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_cri_con_shared_o_status <= 3'd0;
	monroe_ionphoton_cri_con_shared_o_buffer_space_valid <= 1'd0;
	monroe_ionphoton_cri_con_shared_o_buffer_space <= 16'd0;
	monroe_ionphoton_cri_con_shared_i_data <= 32'd0;
	monroe_ionphoton_cri_con_shared_i_timestamp <= 64'd0;
	monroe_ionphoton_cri_con_shared_i_status <= 4'd0;
	case (monroe_ionphoton_cri_con_selected)
		1'd0: begin
			monroe_ionphoton_cri_con_shared_o_status <= monroe_ionphoton_rtio_core_cri_o_status;
			monroe_ionphoton_cri_con_shared_o_buffer_space_valid <= monroe_ionphoton_rtio_core_cri_o_buffer_space_valid;
			monroe_ionphoton_cri_con_shared_o_buffer_space <= monroe_ionphoton_rtio_core_cri_o_buffer_space;
			monroe_ionphoton_cri_con_shared_i_data <= monroe_ionphoton_rtio_core_cri_i_data;
			monroe_ionphoton_cri_con_shared_i_timestamp <= monroe_ionphoton_rtio_core_cri_i_timestamp;
			monroe_ionphoton_cri_con_shared_i_status <= monroe_ionphoton_rtio_core_cri_i_status;
		end
	endcase
// synthesis translate_off
	dummy_d_149 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_r = monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_w[1:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_re = ((((monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank2_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack)) & monroe_ionphoton_monroe_ionphoton_csrbank2_bus_we) & (monroe_ionphoton_monroe_ionphoton_csrbank2_bus_adr[0] == 1'd0));
assign monroe_ionphoton_cri_con_storage = monroe_ionphoton_cri_con_storage_full[1:0];
assign monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_w = monroe_ionphoton_cri_con_storage_full[1:0];
assign monroe_ionphoton_mon_bussynchronizer0_i = inout_8x0_serdes_i0[7];
assign monroe_ionphoton_mon_bussynchronizer1_i = inout_8x0_serdes_oe;
assign monroe_ionphoton_mon_bussynchronizer2_i = inout_8x1_serdes_i0[7];
assign monroe_ionphoton_mon_bussynchronizer3_i = inout_8x1_serdes_oe;
assign monroe_ionphoton_mon_bussynchronizer4_i = inout_8x2_serdes_i0[7];
assign monroe_ionphoton_mon_bussynchronizer5_i = inout_8x2_serdes_oe;
assign monroe_ionphoton_mon_bussynchronizer6_i = inout_8x3_serdes_i0[7];
assign monroe_ionphoton_mon_bussynchronizer7_i = inout_8x3_serdes_oe;
assign monroe_ionphoton_mon_bussynchronizer8_i = output_8x0_o[7];
assign monroe_ionphoton_mon_bussynchronizer9_i = output_8x1_o[7];
assign monroe_ionphoton_mon_bussynchronizer10_i = output_8x2_o[7];
assign monroe_ionphoton_mon_bussynchronizer11_i = output_8x3_o[7];
assign monroe_ionphoton_mon_bussynchronizer12_i = output_8x4_o[7];
assign monroe_ionphoton_mon_bussynchronizer13_i = output_8x5_o[7];
assign monroe_ionphoton_mon_bussynchronizer14_i = output_8x6_o[7];
assign monroe_ionphoton_mon_bussynchronizer15_i = output_8x7_o[7];
assign monroe_ionphoton_mon_bussynchronizer16_i = output_8x8_o[7];
assign monroe_ionphoton_mon_bussynchronizer17_i = output_8x9_o[7];
assign monroe_ionphoton_mon_bussynchronizer18_i = output_8x10_o[7];
assign monroe_ionphoton_mon_bussynchronizer19_i = output_8x11_o[7];
assign monroe_ionphoton_mon_bussynchronizer20_i = output_8x12_o[7];
assign monroe_ionphoton_mon_bussynchronizer21_i = output_8x13_o[7];
assign monroe_ionphoton_mon_bussynchronizer22_i = output_8x14_o[7];
assign monroe_ionphoton_mon_bussynchronizer23_i = output_8x15_o[7];
assign monroe_ionphoton_mon_bussynchronizer24_i = output_8x16_o[7];
assign monroe_ionphoton_mon_bussynchronizer25_i = output_8x17_o[7];
assign monroe_ionphoton_mon_bussynchronizer26_i = output_8x18_o[7];
assign monroe_ionphoton_mon_bussynchronizer27_i = output_8x19_o[7];
assign monroe_ionphoton_mon_bussynchronizer28_i = output_8x20_o[7];
assign monroe_ionphoton_mon_bussynchronizer29_i = output_8x21_o[7];
assign monroe_ionphoton_mon_bussynchronizer30_i = output_8x22_o[7];
assign monroe_ionphoton_mon_bussynchronizer31_i = output_8x23_o[7];
assign monroe_ionphoton_mon_bussynchronizer32_i = output_8x24_o[7];
assign monroe_ionphoton_mon_bussynchronizer33_i = output_8x25_o[7];
assign monroe_ionphoton_mon_bussynchronizer34_i = output_8x26_o[7];
assign monroe_ionphoton_mon_bussynchronizer35_i = output0_pad_o;
assign monroe_ionphoton_mon_bussynchronizer36_i = output1_pad_o;
assign monroe_ionphoton_inj_value_w = comb_rhs_array_muxed16;
assign monroe_ionphoton_rtio_analyzer_fifo_sink_stb = monroe_ionphoton_rtio_analyzer_message_encoder_source_stb;
assign monroe_ionphoton_rtio_analyzer_message_encoder_source_ack = monroe_ionphoton_rtio_analyzer_fifo_sink_ack;
assign monroe_ionphoton_rtio_analyzer_fifo_sink_eop = monroe_ionphoton_rtio_analyzer_message_encoder_source_eop;
assign monroe_ionphoton_rtio_analyzer_fifo_sink_payload_data = monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data;
assign monroe_ionphoton_rtio_analyzer_converter_sink_stb = monroe_ionphoton_rtio_analyzer_fifo_source_stb;
assign monroe_ionphoton_rtio_analyzer_fifo_source_ack = monroe_ionphoton_rtio_analyzer_converter_sink_ack;
assign monroe_ionphoton_rtio_analyzer_converter_sink_eop = monroe_ionphoton_rtio_analyzer_fifo_source_eop;
assign monroe_ionphoton_rtio_analyzer_converter_sink_payload_data = monroe_ionphoton_rtio_analyzer_fifo_source_payload_data;
assign monroe_ionphoton_rtio_analyzer_dma_sink_stb = monroe_ionphoton_rtio_analyzer_converter_source_stb;
assign monroe_ionphoton_rtio_analyzer_converter_source_ack = monroe_ionphoton_rtio_analyzer_dma_sink_ack;
assign monroe_ionphoton_rtio_analyzer_dma_sink_eop = monroe_ionphoton_rtio_analyzer_converter_source_eop;
assign monroe_ionphoton_rtio_analyzer_dma_sink_payload_data = monroe_ionphoton_rtio_analyzer_converter_source_payload_data;
assign monroe_ionphoton_rtio_analyzer_dma_sink_payload_valid_token_count = monroe_ionphoton_rtio_analyzer_converter_source_payload_valid_token_count;

// synthesis translate_off
reg dummy_d_150;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_analyzer_message_encoder_read_done <= 1'd0;
	monroe_ionphoton_rtio_analyzer_message_encoder_read_overflow <= 1'd0;
	if ((monroe_ionphoton_rtio_analyzer_message_encoder_read_wait_event_r & (~monroe_ionphoton_rtio_core_cri_i_status[2]))) begin
		if ((~monroe_ionphoton_rtio_core_cri_i_status[0])) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_read_done <= 1'd1;
		end
		if (monroe_ionphoton_rtio_core_cri_i_status[1]) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_read_overflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_150 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_analyzer_message_encoder_input_output_channel = monroe_ionphoton_rtio_core_cri_chan_sel;
assign monroe_ionphoton_rtio_analyzer_message_encoder_input_output_address_padding = monroe_ionphoton_rtio_core_cri_o_address;
assign monroe_ionphoton_rtio_analyzer_message_encoder_input_output_rtio_counter = monroe_ionphoton_rtio_tsc_full_ts_sys;

// synthesis translate_off
reg dummy_d_151;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_analyzer_message_encoder_input_output_message_type <= 2'd0;
	monroe_ionphoton_rtio_analyzer_message_encoder_input_output_timestamp <= 64'd0;
	monroe_ionphoton_rtio_analyzer_message_encoder_input_output_data <= 64'd0;
	if ((monroe_ionphoton_rtio_core_cri_cmd == 1'd1)) begin
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_message_type <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_timestamp <= monroe_ionphoton_rtio_core_cri_o_timestamp;
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_data <= monroe_ionphoton_rtio_core_cri_o_data;
	end else begin
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_message_type <= 1'd1;
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_timestamp <= monroe_ionphoton_rtio_core_cri_i_timestamp;
		monroe_ionphoton_rtio_analyzer_message_encoder_input_output_data <= monroe_ionphoton_rtio_core_cri_i_data;
	end
// synthesis translate_off
	dummy_d_151 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_analyzer_message_encoder_input_output_stb = ((monroe_ionphoton_rtio_core_cri_cmd == 1'd1) | monroe_ionphoton_rtio_analyzer_message_encoder_read_done);
assign monroe_ionphoton_rtio_analyzer_message_encoder_exception_message_type = 2'd2;
assign monroe_ionphoton_rtio_analyzer_message_encoder_exception_channel = monroe_ionphoton_rtio_core_cri_chan_sel;
assign monroe_ionphoton_rtio_analyzer_message_encoder_exception_rtio_counter = monroe_ionphoton_rtio_tsc_full_ts_sys;

// synthesis translate_off
reg dummy_d_152;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb <= 1'd0;
	monroe_ionphoton_rtio_analyzer_message_encoder_exception_exception_type <= 8'd0;
	if ((monroe_ionphoton_rtio_analyzer_message_encoder_just_written & monroe_ionphoton_rtio_core_cri_o_status[1])) begin
		monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		monroe_ionphoton_rtio_analyzer_message_encoder_exception_exception_type <= 5'd20;
	end
	if (monroe_ionphoton_rtio_analyzer_message_encoder_read_overflow) begin
		monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		monroe_ionphoton_rtio_analyzer_message_encoder_exception_exception_type <= 6'd33;
	end
// synthesis translate_off
	dummy_d_152 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_analyzer_message_encoder_stopped_message_type = 2'd3;
assign monroe_ionphoton_rtio_analyzer_message_encoder_stopped_rtio_counter = monroe_ionphoton_rtio_tsc_full_ts_sys;
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_din = {monroe_ionphoton_rtio_analyzer_fifo_fifo_in_eop, monroe_ionphoton_rtio_analyzer_fifo_fifo_in_payload_data};
assign {monroe_ionphoton_rtio_analyzer_fifo_fifo_out_eop, monroe_ionphoton_rtio_analyzer_fifo_fifo_out_payload_data} = monroe_ionphoton_rtio_analyzer_fifo_syncfifo_dout;
assign monroe_ionphoton_rtio_analyzer_fifo_sink_ack = monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable;
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_we = monroe_ionphoton_rtio_analyzer_fifo_sink_stb;
assign monroe_ionphoton_rtio_analyzer_fifo_fifo_in_eop = monroe_ionphoton_rtio_analyzer_fifo_sink_eop;
assign monroe_ionphoton_rtio_analyzer_fifo_fifo_in_payload_data = monroe_ionphoton_rtio_analyzer_fifo_sink_payload_data;
assign monroe_ionphoton_rtio_analyzer_fifo_source_stb = monroe_ionphoton_rtio_analyzer_fifo_readable;
assign monroe_ionphoton_rtio_analyzer_fifo_source_eop = monroe_ionphoton_rtio_analyzer_fifo_fifo_out_eop;
assign monroe_ionphoton_rtio_analyzer_fifo_source_payload_data = monroe_ionphoton_rtio_analyzer_fifo_fifo_out_payload_data;
assign monroe_ionphoton_rtio_analyzer_fifo_re = monroe_ionphoton_rtio_analyzer_fifo_source_ack;
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_re = (monroe_ionphoton_rtio_analyzer_fifo_syncfifo_readable & ((~monroe_ionphoton_rtio_analyzer_fifo_readable) | monroe_ionphoton_rtio_analyzer_fifo_re));
assign monroe_ionphoton_rtio_analyzer_fifo_level1 = (monroe_ionphoton_rtio_analyzer_fifo_level0 + monroe_ionphoton_rtio_analyzer_fifo_readable);

// synthesis translate_off
reg dummy_d_153;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_analyzer_fifo_wrport_adr <= 7'd0;
	if (monroe_ionphoton_rtio_analyzer_fifo_replace) begin
		monroe_ionphoton_rtio_analyzer_fifo_wrport_adr <= (monroe_ionphoton_rtio_analyzer_fifo_produce - 1'd1);
	end else begin
		monroe_ionphoton_rtio_analyzer_fifo_wrport_adr <= monroe_ionphoton_rtio_analyzer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_153 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_analyzer_fifo_wrport_dat_w = monroe_ionphoton_rtio_analyzer_fifo_syncfifo_din;
assign monroe_ionphoton_rtio_analyzer_fifo_wrport_we = (monroe_ionphoton_rtio_analyzer_fifo_syncfifo_we & (monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable | monroe_ionphoton_rtio_analyzer_fifo_replace));
assign monroe_ionphoton_rtio_analyzer_fifo_do_read = (monroe_ionphoton_rtio_analyzer_fifo_syncfifo_readable & monroe_ionphoton_rtio_analyzer_fifo_syncfifo_re);
assign monroe_ionphoton_rtio_analyzer_fifo_rdport_adr = monroe_ionphoton_rtio_analyzer_fifo_consume;
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_dout = monroe_ionphoton_rtio_analyzer_fifo_rdport_dat_r;
assign monroe_ionphoton_rtio_analyzer_fifo_rdport_re = monroe_ionphoton_rtio_analyzer_fifo_do_read;
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable = (monroe_ionphoton_rtio_analyzer_fifo_level0 != 8'd128);
assign monroe_ionphoton_rtio_analyzer_fifo_syncfifo_readable = (monroe_ionphoton_rtio_analyzer_fifo_level0 != 1'd0);
assign monroe_ionphoton_rtio_analyzer_converter_last = (monroe_ionphoton_rtio_analyzer_converter_mux == 1'd1);
assign monroe_ionphoton_rtio_analyzer_converter_source_stb = monroe_ionphoton_rtio_analyzer_converter_sink_stb;
assign monroe_ionphoton_rtio_analyzer_converter_source_eop = (monroe_ionphoton_rtio_analyzer_converter_sink_eop & monroe_ionphoton_rtio_analyzer_converter_last);
assign monroe_ionphoton_rtio_analyzer_converter_sink_ack = (monroe_ionphoton_rtio_analyzer_converter_last & monroe_ionphoton_rtio_analyzer_converter_source_ack);

// synthesis translate_off
reg dummy_d_154;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_rtio_analyzer_converter_source_payload_data <= 128'd0;
	case (monroe_ionphoton_rtio_analyzer_converter_mux)
		1'd0: begin
			monroe_ionphoton_rtio_analyzer_converter_source_payload_data <= monroe_ionphoton_rtio_analyzer_converter_sink_payload_data[255:128];
		end
		default: begin
			monroe_ionphoton_rtio_analyzer_converter_source_payload_data <= monroe_ionphoton_rtio_analyzer_converter_sink_payload_data[127:0];
		end
	endcase
// synthesis translate_off
	dummy_d_154 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_rtio_analyzer_converter_source_payload_valid_token_count = monroe_ionphoton_rtio_analyzer_converter_last;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_cyc = monroe_ionphoton_rtio_analyzer_dma_sink_stb;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_stb = monroe_ionphoton_rtio_analyzer_dma_sink_stb;
assign monroe_ionphoton_rtio_analyzer_dma_sink_ack = monroe_ionphoton_monroe_ionphoton_interface1_bus_ack;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_we = 1'd1;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_dat_w = monroe_ionphoton_rtio_analyzer_dma_sink_payload_data;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_sel = 16'd65535;
assign monroe_ionphoton_rtio_analyzer_dma_status = (monroe_ionphoton_rtio_analyzer_dma_message_count <<< 3'd5);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr = comb_rhs_array_muxed54;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_w = comb_rhs_array_muxed55;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_sel = comb_rhs_array_muxed56;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cyc = comb_rhs_array_muxed57;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_stb = comb_rhs_array_muxed58;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_we = comb_rhs_array_muxed59;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_cti = comb_rhs_array_muxed60;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_bte = comb_rhs_array_muxed61;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r;
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_ack = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack & (sdram_cpulevel_arbiter_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_ack = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_ack & (sdram_cpulevel_arbiter_grant == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_err = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_err & (sdram_cpulevel_arbiter_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_err = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_err & (sdram_cpulevel_arbiter_grant == 1'd1));
assign sdram_cpulevel_arbiter_request = {(monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cyc & (~monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_ack)), (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cyc & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_ack))};
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_adr = comb_rhs_array_muxed62;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_w = comb_rhs_array_muxed63;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_sel = comb_rhs_array_muxed64;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_cyc = comb_rhs_array_muxed65;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_stb = comb_rhs_array_muxed66;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_we = comb_rhs_array_muxed67;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_cti = comb_rhs_array_muxed68;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_bte = comb_rhs_array_muxed69;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_r;
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_r;
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_dat_r = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_ack = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack & (sdram_native_arbiter_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_ack = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack & (sdram_native_arbiter_grant == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_ack = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_ack & (sdram_native_arbiter_grant == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_err = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_err & (sdram_native_arbiter_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_interface0_bus_err = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_err & (sdram_native_arbiter_grant == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_interface1_bus_err = (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bus_err & (sdram_native_arbiter_grant == 2'd2));
assign sdram_native_arbiter_request = {(monroe_ionphoton_monroe_ionphoton_interface1_bus_cyc & (~monroe_ionphoton_monroe_ionphoton_interface1_bus_ack)), (monroe_ionphoton_monroe_ionphoton_interface0_bus_cyc & (~monroe_ionphoton_monroe_ionphoton_interface0_bus_ack)), (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_ack))};
assign monroe_ionphoton_shared_adr = comb_rhs_array_muxed70;
assign monroe_ionphoton_shared_dat_w = comb_rhs_array_muxed71;
assign monroe_ionphoton_shared_sel = comb_rhs_array_muxed72;
assign monroe_ionphoton_shared_cyc = comb_rhs_array_muxed73;
assign monroe_ionphoton_shared_stb = comb_rhs_array_muxed74;
assign monroe_ionphoton_shared_we = comb_rhs_array_muxed75;
assign monroe_ionphoton_shared_cti = comb_rhs_array_muxed76;
assign monroe_ionphoton_shared_bte = comb_rhs_array_muxed77;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_r = monroe_ionphoton_shared_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_r = monroe_ionphoton_shared_dat_r;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_ack = (monroe_ionphoton_shared_ack & (monroe_ionphoton_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_ack = (monroe_ionphoton_shared_ack & (monroe_ionphoton_grant == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_err = (monroe_ionphoton_shared_err & (monroe_ionphoton_grant == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_err = (monroe_ionphoton_shared_err & (monroe_ionphoton_grant == 1'd1));
assign monroe_ionphoton_request = {(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cyc & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_ack)), (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cyc & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_ack))};

// synthesis translate_off
reg dummy_d_155;
// synthesis translate_on
always @(*) begin
	monroe_ionphoton_slave_sel <= 6'd0;
	monroe_ionphoton_slave_sel[0] <= (((1'd1 & (~monroe_ionphoton_shared_adr[27])) & (~monroe_ionphoton_shared_adr[28])) & monroe_ionphoton_shared_adr[26]);
	monroe_ionphoton_slave_sel[1] <= (((1'd1 & (~monroe_ionphoton_shared_adr[26])) & monroe_ionphoton_shared_adr[27]) & monroe_ionphoton_shared_adr[28]);
	monroe_ionphoton_slave_sel[2] <= ((1'd1 & (~monroe_ionphoton_shared_adr[27])) & monroe_ionphoton_shared_adr[28]);
	monroe_ionphoton_slave_sel[3] <= (((1'd1 & (~monroe_ionphoton_shared_adr[26])) & (~monroe_ionphoton_shared_adr[27])) & (~monroe_ionphoton_shared_adr[28]));
	monroe_ionphoton_slave_sel[4] <= ((1'd1 & (~monroe_ionphoton_shared_adr[28])) & monroe_ionphoton_shared_adr[27]);
	monroe_ionphoton_slave_sel[5] <= (((1'd1 & monroe_ionphoton_shared_adr[26]) & monroe_ionphoton_shared_adr[27]) & monroe_ionphoton_shared_adr[28]);
// synthesis translate_off
	dummy_d_155 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_bus_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_bus_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_bus_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_bus_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_bus_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_bus_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_bus_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_adr = monroe_ionphoton_shared_adr;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_w = monroe_ionphoton_shared_dat_w;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_sel = monroe_ionphoton_shared_sel;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_stb = monroe_ionphoton_shared_stb;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_we = monroe_ionphoton_shared_we;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_cti = monroe_ionphoton_shared_cti;
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_bte = monroe_ionphoton_shared_bte;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[0]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[1]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[2]);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[3]);
assign monroe_ionphoton_monroe_ionphoton_bus_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[4]);
assign monroe_ionphoton_monroe_ionphoton_mailbox_i1_cyc = (monroe_ionphoton_shared_cyc & monroe_ionphoton_slave_sel[5]);
assign monroe_ionphoton_shared_ack = (((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_ack) | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_ack) | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_ack) | monroe_ionphoton_monroe_ionphoton_bus_ack) | monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack);
assign monroe_ionphoton_shared_err = (((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_err | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_err) | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_err) | monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_err) | monroe_ionphoton_monroe_ionphoton_bus_err) | monroe_ionphoton_monroe_ionphoton_mailbox_i1_err);
assign monroe_ionphoton_shared_dat_r = (((((({32{monroe_ionphoton_slave_sel_r[0]}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_dat_r) | ({32{monroe_ionphoton_slave_sel_r[1]}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_r)) | ({32{monroe_ionphoton_slave_sel_r[2]}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_r)) | ({32{monroe_ionphoton_slave_sel_r[3]}} & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_dat_r)) | ({32{monroe_ionphoton_slave_sel_r[4]}} & monroe_ionphoton_monroe_ionphoton_bus_dat_r)) | ({32{monroe_ionphoton_slave_sel_r[5]}} & monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_r));
assign monroe_ionphoton_csrbank0_sel = (monroe_ionphoton_interface0_bank_bus_adr[13:9] == 3'd7);
assign monroe_ionphoton_csrbank0_dly_sel0_r = monroe_ionphoton_interface0_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank0_dly_sel0_re = ((monroe_ionphoton_csrbank0_sel & monroe_ionphoton_interface0_bank_bus_we) & (monroe_ionphoton_interface0_bank_bus_adr[1:0] == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_r = monroe_ionphoton_interface0_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re = ((monroe_ionphoton_csrbank0_sel & monroe_ionphoton_interface0_bank_bus_we) & (monroe_ionphoton_interface0_bank_bus_adr[1:0] == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_r = monroe_ionphoton_interface0_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re = ((monroe_ionphoton_csrbank0_sel & monroe_ionphoton_interface0_bank_bus_we) & (monroe_ionphoton_interface0_bank_bus_adr[1:0] == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_r = monroe_ionphoton_interface0_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re = ((monroe_ionphoton_csrbank0_sel & monroe_ionphoton_interface0_bank_bus_we) & (monroe_ionphoton_interface0_bank_bus_adr[1:0] == 2'd3));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage_full[1:0];
assign monroe_ionphoton_csrbank0_dly_sel0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage_full[1:0];
assign monroe_ionphoton_csrbank1_sel = (monroe_ionphoton_interface1_bank_bus_adr[13:9] == 3'd5);
assign monroe_ionphoton_csrbank1_control0_r = monroe_ionphoton_interface1_bank_bus_dat_w[3:0];
assign monroe_ionphoton_csrbank1_control0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 1'd0));
assign monroe_ionphoton_csrbank1_pi0_command0_r = monroe_ionphoton_interface1_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank1_pi0_command0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 1'd1));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_r = monroe_ionphoton_interface1_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 2'd2));
assign monroe_ionphoton_csrbank1_pi0_address1_r = monroe_ionphoton_interface1_bank_bus_dat_w[6:0];
assign monroe_ionphoton_csrbank1_pi0_address1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 2'd3));
assign monroe_ionphoton_csrbank1_pi0_address0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_address0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 3'd4));
assign monroe_ionphoton_csrbank1_pi0_baddress0_r = monroe_ionphoton_interface1_bank_bus_dat_w[2:0];
assign monroe_ionphoton_csrbank1_pi0_baddress0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 3'd5));
assign monroe_ionphoton_csrbank1_pi0_wrdata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_wrdata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 3'd6));
assign monroe_ionphoton_csrbank1_pi0_wrdata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_wrdata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 3'd7));
assign monroe_ionphoton_csrbank1_pi0_wrdata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_wrdata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd8));
assign monroe_ionphoton_csrbank1_pi0_wrdata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_wrdata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd9));
assign monroe_ionphoton_csrbank1_pi0_rddata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_rddata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd10));
assign monroe_ionphoton_csrbank1_pi0_rddata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_rddata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd11));
assign monroe_ionphoton_csrbank1_pi0_rddata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_rddata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd12));
assign monroe_ionphoton_csrbank1_pi0_rddata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi0_rddata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd13));
assign monroe_ionphoton_csrbank1_pi1_command0_r = monroe_ionphoton_interface1_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank1_pi1_command0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd14));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_r = monroe_ionphoton_interface1_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 4'd15));
assign monroe_ionphoton_csrbank1_pi1_address1_r = monroe_ionphoton_interface1_bank_bus_dat_w[6:0];
assign monroe_ionphoton_csrbank1_pi1_address1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd16));
assign monroe_ionphoton_csrbank1_pi1_address0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_address0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd17));
assign monroe_ionphoton_csrbank1_pi1_baddress0_r = monroe_ionphoton_interface1_bank_bus_dat_w[2:0];
assign monroe_ionphoton_csrbank1_pi1_baddress0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd18));
assign monroe_ionphoton_csrbank1_pi1_wrdata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_wrdata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd19));
assign monroe_ionphoton_csrbank1_pi1_wrdata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_wrdata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd20));
assign monroe_ionphoton_csrbank1_pi1_wrdata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_wrdata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd21));
assign monroe_ionphoton_csrbank1_pi1_wrdata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_wrdata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd22));
assign monroe_ionphoton_csrbank1_pi1_rddata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_rddata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd23));
assign monroe_ionphoton_csrbank1_pi1_rddata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_rddata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd24));
assign monroe_ionphoton_csrbank1_pi1_rddata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_rddata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd25));
assign monroe_ionphoton_csrbank1_pi1_rddata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi1_rddata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd26));
assign monroe_ionphoton_csrbank1_pi2_command0_r = monroe_ionphoton_interface1_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank1_pi2_command0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd27));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_r = monroe_ionphoton_interface1_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd28));
assign monroe_ionphoton_csrbank1_pi2_address1_r = monroe_ionphoton_interface1_bank_bus_dat_w[6:0];
assign monroe_ionphoton_csrbank1_pi2_address1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd29));
assign monroe_ionphoton_csrbank1_pi2_address0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_address0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd30));
assign monroe_ionphoton_csrbank1_pi2_baddress0_r = monroe_ionphoton_interface1_bank_bus_dat_w[2:0];
assign monroe_ionphoton_csrbank1_pi2_baddress0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 5'd31));
assign monroe_ionphoton_csrbank1_pi2_wrdata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_wrdata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd32));
assign monroe_ionphoton_csrbank1_pi2_wrdata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_wrdata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd33));
assign monroe_ionphoton_csrbank1_pi2_wrdata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_wrdata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd34));
assign monroe_ionphoton_csrbank1_pi2_wrdata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_wrdata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd35));
assign monroe_ionphoton_csrbank1_pi2_rddata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_rddata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd36));
assign monroe_ionphoton_csrbank1_pi2_rddata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_rddata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd37));
assign monroe_ionphoton_csrbank1_pi2_rddata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_rddata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd38));
assign monroe_ionphoton_csrbank1_pi2_rddata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi2_rddata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd39));
assign monroe_ionphoton_csrbank1_pi3_command0_r = monroe_ionphoton_interface1_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank1_pi3_command0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd40));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_r = monroe_ionphoton_interface1_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd41));
assign monroe_ionphoton_csrbank1_pi3_address1_r = monroe_ionphoton_interface1_bank_bus_dat_w[6:0];
assign monroe_ionphoton_csrbank1_pi3_address1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd42));
assign monroe_ionphoton_csrbank1_pi3_address0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_address0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd43));
assign monroe_ionphoton_csrbank1_pi3_baddress0_r = monroe_ionphoton_interface1_bank_bus_dat_w[2:0];
assign monroe_ionphoton_csrbank1_pi3_baddress0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd44));
assign monroe_ionphoton_csrbank1_pi3_wrdata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_wrdata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd45));
assign monroe_ionphoton_csrbank1_pi3_wrdata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_wrdata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd46));
assign monroe_ionphoton_csrbank1_pi3_wrdata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_wrdata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd47));
assign monroe_ionphoton_csrbank1_pi3_wrdata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_wrdata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd48));
assign monroe_ionphoton_csrbank1_pi3_rddata3_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_rddata3_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd49));
assign monroe_ionphoton_csrbank1_pi3_rddata2_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_rddata2_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd50));
assign monroe_ionphoton_csrbank1_pi3_rddata1_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_rddata1_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd51));
assign monroe_ionphoton_csrbank1_pi3_rddata0_r = monroe_ionphoton_interface1_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank1_pi3_rddata0_re = ((monroe_ionphoton_csrbank1_sel & monroe_ionphoton_interface1_bank_bus_we) & (monroe_ionphoton_interface1_bank_bus_adr[5:0] == 6'd52));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage_full[3:0];
assign monroe_ionphoton_csrbank1_control0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage_full[3:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage_full[5:0];
assign monroe_ionphoton_csrbank1_pi0_command0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage_full[5:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full[14:0];
assign monroe_ionphoton_csrbank1_pi0_address1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full[14:8];
assign monroe_ionphoton_csrbank1_pi0_address0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage_full[2:0];
assign monroe_ionphoton_csrbank1_pi0_baddress0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage_full[2:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[31:0];
assign monroe_ionphoton_csrbank1_pi0_wrdata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[31:24];
assign monroe_ionphoton_csrbank1_pi0_wrdata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[23:16];
assign monroe_ionphoton_csrbank1_pi0_wrdata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[15:8];
assign monroe_ionphoton_csrbank1_pi0_wrdata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[7:0];
assign monroe_ionphoton_csrbank1_pi0_rddata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status[31:24];
assign monroe_ionphoton_csrbank1_pi0_rddata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status[23:16];
assign monroe_ionphoton_csrbank1_pi0_rddata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status[15:8];
assign monroe_ionphoton_csrbank1_pi0_rddata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage_full[5:0];
assign monroe_ionphoton_csrbank1_pi1_command0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage_full[5:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full[14:0];
assign monroe_ionphoton_csrbank1_pi1_address1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full[14:8];
assign monroe_ionphoton_csrbank1_pi1_address0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage_full[2:0];
assign monroe_ionphoton_csrbank1_pi1_baddress0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage_full[2:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[31:0];
assign monroe_ionphoton_csrbank1_pi1_wrdata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[31:24];
assign monroe_ionphoton_csrbank1_pi1_wrdata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[23:16];
assign monroe_ionphoton_csrbank1_pi1_wrdata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[15:8];
assign monroe_ionphoton_csrbank1_pi1_wrdata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[7:0];
assign monroe_ionphoton_csrbank1_pi1_rddata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status[31:24];
assign monroe_ionphoton_csrbank1_pi1_rddata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status[23:16];
assign monroe_ionphoton_csrbank1_pi1_rddata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status[15:8];
assign monroe_ionphoton_csrbank1_pi1_rddata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage_full[5:0];
assign monroe_ionphoton_csrbank1_pi2_command0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage_full[5:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full[14:0];
assign monroe_ionphoton_csrbank1_pi2_address1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full[14:8];
assign monroe_ionphoton_csrbank1_pi2_address0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage_full[2:0];
assign monroe_ionphoton_csrbank1_pi2_baddress0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage_full[2:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[31:0];
assign monroe_ionphoton_csrbank1_pi2_wrdata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[31:24];
assign monroe_ionphoton_csrbank1_pi2_wrdata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[23:16];
assign monroe_ionphoton_csrbank1_pi2_wrdata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[15:8];
assign monroe_ionphoton_csrbank1_pi2_wrdata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[7:0];
assign monroe_ionphoton_csrbank1_pi2_rddata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status[31:24];
assign monroe_ionphoton_csrbank1_pi2_rddata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status[23:16];
assign monroe_ionphoton_csrbank1_pi2_rddata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status[15:8];
assign monroe_ionphoton_csrbank1_pi2_rddata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage_full[5:0];
assign monroe_ionphoton_csrbank1_pi3_command0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage_full[5:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full[14:0];
assign monroe_ionphoton_csrbank1_pi3_address1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full[14:8];
assign monroe_ionphoton_csrbank1_pi3_address0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage_full[2:0];
assign monroe_ionphoton_csrbank1_pi3_baddress0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage_full[2:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[31:0];
assign monroe_ionphoton_csrbank1_pi3_wrdata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[31:24];
assign monroe_ionphoton_csrbank1_pi3_wrdata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[23:16];
assign monroe_ionphoton_csrbank1_pi3_wrdata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[15:8];
assign monroe_ionphoton_csrbank1_pi3_wrdata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[7:0];
assign monroe_ionphoton_csrbank1_pi3_rddata3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status[31:24];
assign monroe_ionphoton_csrbank1_pi3_rddata2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status[23:16];
assign monroe_ionphoton_csrbank1_pi3_rddata1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status[15:8];
assign monroe_ionphoton_csrbank1_pi3_rddata0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status[7:0];
assign monroe_ionphoton_csrbank2_sel = (monroe_ionphoton_interface2_bank_bus_adr[13:9] == 4'd10);
assign monroe_ionphoton_csrbank2_sram_writer_slot_r = monroe_ionphoton_interface2_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank2_sram_writer_slot_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 1'd0));
assign monroe_ionphoton_csrbank2_sram_writer_length3_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_length3_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 1'd1));
assign monroe_ionphoton_csrbank2_sram_writer_length2_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_length2_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 2'd2));
assign monroe_ionphoton_csrbank2_sram_writer_length1_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_length1_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 2'd3));
assign monroe_ionphoton_csrbank2_sram_writer_length0_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_length0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 3'd4));
assign monroe_ionphoton_csrbank2_sram_writer_errors3_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_errors3_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 3'd5));
assign monroe_ionphoton_csrbank2_sram_writer_errors2_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_errors2_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 3'd6));
assign monroe_ionphoton_csrbank2_sram_writer_errors1_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_errors1_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 3'd7));
assign monroe_ionphoton_csrbank2_sram_writer_errors0_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_errors0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd8));
assign monroe_ionphoton_monroe_ionphoton_writer_status_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_writer_status_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd9));
assign monroe_ionphoton_monroe_ionphoton_writer_pending_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_writer_pending_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd10));
assign monroe_ionphoton_csrbank2_sram_writer_ev_enable0_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank2_sram_writer_ev_enable0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd11));
assign monroe_ionphoton_monroe_ionphoton_reader_start_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_reader_start_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd12));
assign monroe_ionphoton_csrbank2_sram_reader_ready_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank2_sram_reader_ready_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd13));
assign monroe_ionphoton_csrbank2_sram_reader_slot0_r = monroe_ionphoton_interface2_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank2_sram_reader_slot0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd14));
assign monroe_ionphoton_csrbank2_sram_reader_length1_r = monroe_ionphoton_interface2_bank_bus_dat_w[2:0];
assign monroe_ionphoton_csrbank2_sram_reader_length1_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 4'd15));
assign monroe_ionphoton_csrbank2_sram_reader_length0_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_sram_reader_length0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd16));
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd17));
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd18));
assign monroe_ionphoton_csrbank2_sram_reader_ev_enable0_r = monroe_ionphoton_interface2_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank2_sram_reader_ev_enable0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd19));
assign monroe_ionphoton_csrbank2_preamble_errors3_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_preamble_errors3_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd20));
assign monroe_ionphoton_csrbank2_preamble_errors2_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_preamble_errors2_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd21));
assign monroe_ionphoton_csrbank2_preamble_errors1_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_preamble_errors1_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd22));
assign monroe_ionphoton_csrbank2_preamble_errors0_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_preamble_errors0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd23));
assign monroe_ionphoton_csrbank2_crc_errors3_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_crc_errors3_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd24));
assign monroe_ionphoton_csrbank2_crc_errors2_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_crc_errors2_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd25));
assign monroe_ionphoton_csrbank2_crc_errors1_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_crc_errors1_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd26));
assign monroe_ionphoton_csrbank2_crc_errors0_r = monroe_ionphoton_interface2_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank2_crc_errors0_re = ((monroe_ionphoton_csrbank2_sel & monroe_ionphoton_interface2_bank_bus_we) & (monroe_ionphoton_interface2_bank_bus_adr[4:0] == 5'd27));
assign monroe_ionphoton_csrbank2_sram_writer_slot_w = monroe_ionphoton_monroe_ionphoton_writer_slot_status[1:0];
assign monroe_ionphoton_csrbank2_sram_writer_length3_w = monroe_ionphoton_monroe_ionphoton_writer_length_status[31:24];
assign monroe_ionphoton_csrbank2_sram_writer_length2_w = monroe_ionphoton_monroe_ionphoton_writer_length_status[23:16];
assign monroe_ionphoton_csrbank2_sram_writer_length1_w = monroe_ionphoton_monroe_ionphoton_writer_length_status[15:8];
assign monroe_ionphoton_csrbank2_sram_writer_length0_w = monroe_ionphoton_monroe_ionphoton_writer_length_status[7:0];
assign monroe_ionphoton_csrbank2_sram_writer_errors3_w = monroe_ionphoton_monroe_ionphoton_writer_errors_status[31:24];
assign monroe_ionphoton_csrbank2_sram_writer_errors2_w = monroe_ionphoton_monroe_ionphoton_writer_errors_status[23:16];
assign monroe_ionphoton_csrbank2_sram_writer_errors1_w = monroe_ionphoton_monroe_ionphoton_writer_errors_status[15:8];
assign monroe_ionphoton_csrbank2_sram_writer_errors0_w = monroe_ionphoton_monroe_ionphoton_writer_errors_status[7:0];
assign monroe_ionphoton_monroe_ionphoton_writer_storage = monroe_ionphoton_monroe_ionphoton_writer_storage_full;
assign monroe_ionphoton_csrbank2_sram_writer_ev_enable0_w = monroe_ionphoton_monroe_ionphoton_writer_storage_full;
assign monroe_ionphoton_csrbank2_sram_reader_ready_w = monroe_ionphoton_monroe_ionphoton_reader_ready_status;
assign monroe_ionphoton_monroe_ionphoton_reader_slot_storage = monroe_ionphoton_monroe_ionphoton_reader_slot_storage_full[1:0];
assign monroe_ionphoton_csrbank2_sram_reader_slot0_w = monroe_ionphoton_monroe_ionphoton_reader_slot_storage_full[1:0];
assign monroe_ionphoton_monroe_ionphoton_reader_length_storage = monroe_ionphoton_monroe_ionphoton_reader_length_storage_full[10:0];
assign monroe_ionphoton_csrbank2_sram_reader_length1_w = monroe_ionphoton_monroe_ionphoton_reader_length_storage_full[10:8];
assign monroe_ionphoton_csrbank2_sram_reader_length0_w = monroe_ionphoton_monroe_ionphoton_reader_length_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage = monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage_full;
assign monroe_ionphoton_csrbank2_sram_reader_ev_enable0_w = monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage_full;
assign monroe_ionphoton_csrbank2_preamble_errors3_w = monroe_ionphoton_monroe_ionphoton_preamble_errors_status[31:24];
assign monroe_ionphoton_csrbank2_preamble_errors2_w = monroe_ionphoton_monroe_ionphoton_preamble_errors_status[23:16];
assign monroe_ionphoton_csrbank2_preamble_errors1_w = monroe_ionphoton_monroe_ionphoton_preamble_errors_status[15:8];
assign monroe_ionphoton_csrbank2_preamble_errors0_w = monroe_ionphoton_monroe_ionphoton_preamble_errors_status[7:0];
assign monroe_ionphoton_csrbank2_crc_errors3_w = monroe_ionphoton_monroe_ionphoton_crc_errors_status[31:24];
assign monroe_ionphoton_csrbank2_crc_errors2_w = monroe_ionphoton_monroe_ionphoton_crc_errors_status[23:16];
assign monroe_ionphoton_csrbank2_crc_errors1_w = monroe_ionphoton_monroe_ionphoton_crc_errors_status[15:8];
assign monroe_ionphoton_csrbank2_crc_errors0_w = monroe_ionphoton_monroe_ionphoton_crc_errors_status[7:0];
assign monroe_ionphoton_csrbank3_sel = (monroe_ionphoton_interface3_bank_bus_adr[13:9] == 4'd13);
assign monroe_ionphoton_csrbank3_in_r = monroe_ionphoton_interface3_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank3_in_re = ((monroe_ionphoton_csrbank3_sel & monroe_ionphoton_interface3_bank_bus_we) & (monroe_ionphoton_interface3_bank_bus_adr[1:0] == 1'd0));
assign monroe_ionphoton_csrbank3_out0_r = monroe_ionphoton_interface3_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank3_out0_re = ((monroe_ionphoton_csrbank3_sel & monroe_ionphoton_interface3_bank_bus_we) & (monroe_ionphoton_interface3_bank_bus_adr[1:0] == 1'd1));
assign monroe_ionphoton_csrbank3_oe0_r = monroe_ionphoton_interface3_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank3_oe0_re = ((monroe_ionphoton_csrbank3_sel & monroe_ionphoton_interface3_bank_bus_we) & (monroe_ionphoton_interface3_bank_bus_adr[1:0] == 2'd2));
assign monroe_ionphoton_csrbank3_in_w = monroe_ionphoton_i2c_status0[1:0];
assign monroe_ionphoton_i2c_out_storage = monroe_ionphoton_i2c_out_storage_full[1:0];
assign monroe_ionphoton_csrbank3_out0_w = monroe_ionphoton_i2c_out_storage_full[1:0];
assign monroe_ionphoton_i2c_oe_storage = monroe_ionphoton_i2c_oe_storage_full[1:0];
assign monroe_ionphoton_csrbank3_oe0_w = monroe_ionphoton_i2c_oe_storage_full[1:0];
assign monroe_ionphoton_csrbank4_sel = (monroe_ionphoton_interface4_bank_bus_adr[13:9] == 2'd2);
assign monroe_ionphoton_csrbank4_address0_r = monroe_ionphoton_interface4_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank4_address0_re = ((monroe_ionphoton_csrbank4_sel & monroe_ionphoton_interface4_bank_bus_we) & (monroe_ionphoton_interface4_bank_bus_adr[0] == 1'd0));
assign monroe_ionphoton_csrbank4_data_r = monroe_ionphoton_interface4_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank4_data_re = ((monroe_ionphoton_csrbank4_sel & monroe_ionphoton_interface4_bank_bus_we) & (monroe_ionphoton_interface4_bank_bus_adr[0] == 1'd1));
assign monroe_ionphoton_add_identifier_storage = monroe_ionphoton_add_identifier_storage_full[7:0];
assign monroe_ionphoton_csrbank4_address0_w = monroe_ionphoton_add_identifier_storage_full[7:0];
assign monroe_ionphoton_csrbank4_data_w = monroe_ionphoton_add_identifier_status[7:0];
assign monroe_ionphoton_csrbank5_sel = (monroe_ionphoton_interface5_bank_bus_adr[13:9] == 4'd11);
assign monroe_ionphoton_csrbank5_reset0_r = monroe_ionphoton_interface5_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank5_reset0_re = ((monroe_ionphoton_csrbank5_sel & monroe_ionphoton_interface5_bank_bus_we) & (monroe_ionphoton_interface5_bank_bus_adr[0] == 1'd0));
assign monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage = monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage_full;
assign monroe_ionphoton_csrbank5_reset0_w = monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage_full;
assign monroe_ionphoton_csrbank6_sel = (monroe_ionphoton_interface6_bank_bus_adr[13:9] == 4'd12);
assign monroe_ionphoton_csrbank6_out0_r = monroe_ionphoton_interface6_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank6_out0_re = ((monroe_ionphoton_csrbank6_sel & monroe_ionphoton_interface6_bank_bus_we) & (monroe_ionphoton_interface6_bank_bus_adr[0] == 1'd0));
assign monroe_ionphoton_leds_storage = monroe_ionphoton_leds_storage_full;
assign monroe_ionphoton_csrbank6_out0_w = monroe_ionphoton_leds_storage_full;
assign monroe_ionphoton_csrbank7_sel = (monroe_ionphoton_interface7_bank_bus_adr[13:9] == 5'd17);
assign monroe_ionphoton_csrbank7_enable0_r = monroe_ionphoton_interface7_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank7_enable0_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 1'd0));
assign monroe_ionphoton_csrbank7_busy_r = monroe_ionphoton_interface7_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank7_busy_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 1'd1));
assign monroe_ionphoton_csrbank7_message_encoder_overflow_r = monroe_ionphoton_interface7_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank7_message_encoder_overflow_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 2'd2));
assign monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_r = monroe_ionphoton_interface7_bank_bus_dat_w[0];
assign monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 2'd3));
assign monroe_ionphoton_rtio_analyzer_dma_reset_r = monroe_ionphoton_interface7_bank_bus_dat_w[0];
assign monroe_ionphoton_rtio_analyzer_dma_reset_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 3'd4));
assign monroe_ionphoton_csrbank7_dma_base_address4_r = monroe_ionphoton_interface7_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank7_dma_base_address4_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 3'd5));
assign monroe_ionphoton_csrbank7_dma_base_address3_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_base_address3_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 3'd6));
assign monroe_ionphoton_csrbank7_dma_base_address2_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_base_address2_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 3'd7));
assign monroe_ionphoton_csrbank7_dma_base_address1_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_base_address1_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd8));
assign monroe_ionphoton_csrbank7_dma_base_address0_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_base_address0_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd9));
assign monroe_ionphoton_csrbank7_dma_last_address4_r = monroe_ionphoton_interface7_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank7_dma_last_address4_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd10));
assign monroe_ionphoton_csrbank7_dma_last_address3_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_last_address3_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd11));
assign monroe_ionphoton_csrbank7_dma_last_address2_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_last_address2_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd12));
assign monroe_ionphoton_csrbank7_dma_last_address1_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_last_address1_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd13));
assign monroe_ionphoton_csrbank7_dma_last_address0_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_last_address0_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd14));
assign monroe_ionphoton_csrbank7_dma_byte_count7_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count7_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 4'd15));
assign monroe_ionphoton_csrbank7_dma_byte_count6_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count6_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd16));
assign monroe_ionphoton_csrbank7_dma_byte_count5_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count5_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd17));
assign monroe_ionphoton_csrbank7_dma_byte_count4_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count4_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd18));
assign monroe_ionphoton_csrbank7_dma_byte_count3_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count3_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd19));
assign monroe_ionphoton_csrbank7_dma_byte_count2_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count2_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd20));
assign monroe_ionphoton_csrbank7_dma_byte_count1_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count1_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd21));
assign monroe_ionphoton_csrbank7_dma_byte_count0_r = monroe_ionphoton_interface7_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank7_dma_byte_count0_re = ((monroe_ionphoton_csrbank7_sel & monroe_ionphoton_interface7_bank_bus_we) & (monroe_ionphoton_interface7_bank_bus_adr[4:0] == 5'd22));
assign monroe_ionphoton_rtio_analyzer_enable_storage = monroe_ionphoton_rtio_analyzer_enable_storage_full;
assign monroe_ionphoton_csrbank7_enable0_w = monroe_ionphoton_rtio_analyzer_enable_storage_full;
assign monroe_ionphoton_csrbank7_busy_w = monroe_ionphoton_rtio_analyzer_busy_status;
assign monroe_ionphoton_csrbank7_message_encoder_overflow_w = monroe_ionphoton_rtio_analyzer_message_encoder_status;
assign monroe_ionphoton_rtio_analyzer_dma_base_address_storage = monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[33:4];
assign monroe_ionphoton_csrbank7_dma_base_address4_w = monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[33:32];
assign monroe_ionphoton_csrbank7_dma_base_address3_w = monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[31:24];
assign monroe_ionphoton_csrbank7_dma_base_address2_w = monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[23:16];
assign monroe_ionphoton_csrbank7_dma_base_address1_w = monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[15:8];
assign monroe_ionphoton_csrbank7_dma_base_address0_w = {monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[7:4], {4{1'd0}}};
assign monroe_ionphoton_rtio_analyzer_dma_last_address_storage = monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[33:4];
assign monroe_ionphoton_csrbank7_dma_last_address4_w = monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[33:32];
assign monroe_ionphoton_csrbank7_dma_last_address3_w = monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[31:24];
assign monroe_ionphoton_csrbank7_dma_last_address2_w = monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[23:16];
assign monroe_ionphoton_csrbank7_dma_last_address1_w = monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[15:8];
assign monroe_ionphoton_csrbank7_dma_last_address0_w = {monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[7:4], {4{1'd0}}};
assign monroe_ionphoton_csrbank7_dma_byte_count7_w = monroe_ionphoton_rtio_analyzer_dma_status[63:56];
assign monroe_ionphoton_csrbank7_dma_byte_count6_w = monroe_ionphoton_rtio_analyzer_dma_status[55:48];
assign monroe_ionphoton_csrbank7_dma_byte_count5_w = monroe_ionphoton_rtio_analyzer_dma_status[47:40];
assign monroe_ionphoton_csrbank7_dma_byte_count4_w = monroe_ionphoton_rtio_analyzer_dma_status[39:32];
assign monroe_ionphoton_csrbank7_dma_byte_count3_w = monroe_ionphoton_rtio_analyzer_dma_status[31:24];
assign monroe_ionphoton_csrbank7_dma_byte_count2_w = monroe_ionphoton_rtio_analyzer_dma_status[23:16];
assign monroe_ionphoton_csrbank7_dma_byte_count1_w = monroe_ionphoton_rtio_analyzer_dma_status[15:8];
assign monroe_ionphoton_csrbank7_dma_byte_count0_w = monroe_ionphoton_rtio_analyzer_dma_status[7:0];
assign monroe_ionphoton_csrbank8_sel = (monroe_ionphoton_interface8_bank_bus_adr[13:9] == 4'd15);
assign monroe_ionphoton_rtio_core_reset_r = monroe_ionphoton_interface8_bank_bus_dat_w[0];
assign monroe_ionphoton_rtio_core_reset_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 1'd0));
assign monroe_ionphoton_rtio_core_reset_phy_r = monroe_ionphoton_interface8_bank_bus_dat_w[0];
assign monroe_ionphoton_rtio_core_reset_phy_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 1'd1));
assign monroe_ionphoton_rtio_core_async_error_r = monroe_ionphoton_interface8_bank_bus_dat_w[2:0];
assign monroe_ionphoton_rtio_core_async_error_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 2'd2));
assign monroe_ionphoton_csrbank8_collision_channel1_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_collision_channel1_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 2'd3));
assign monroe_ionphoton_csrbank8_collision_channel0_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_collision_channel0_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 3'd4));
assign monroe_ionphoton_csrbank8_busy_channel1_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_busy_channel1_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 3'd5));
assign monroe_ionphoton_csrbank8_busy_channel0_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_busy_channel0_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 3'd6));
assign monroe_ionphoton_csrbank8_sequence_error_channel1_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_sequence_error_channel1_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 3'd7));
assign monroe_ionphoton_csrbank8_sequence_error_channel0_r = monroe_ionphoton_interface8_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank8_sequence_error_channel0_re = ((monroe_ionphoton_csrbank8_sel & monroe_ionphoton_interface8_bank_bus_we) & (monroe_ionphoton_interface8_bank_bus_adr[3:0] == 4'd8));
assign monroe_ionphoton_csrbank8_collision_channel1_w = monroe_ionphoton_rtio_core_collision_channel_status[15:8];
assign monroe_ionphoton_csrbank8_collision_channel0_w = monroe_ionphoton_rtio_core_collision_channel_status[7:0];
assign monroe_ionphoton_csrbank8_busy_channel1_w = monroe_ionphoton_rtio_core_busy_channel_status[15:8];
assign monroe_ionphoton_csrbank8_busy_channel0_w = monroe_ionphoton_rtio_core_busy_channel_status[7:0];
assign monroe_ionphoton_csrbank8_sequence_error_channel1_w = monroe_ionphoton_rtio_core_sequence_error_channel_status[15:8];
assign monroe_ionphoton_csrbank8_sequence_error_channel0_w = monroe_ionphoton_rtio_core_sequence_error_channel_status[7:0];
assign monroe_ionphoton_csrbank9_sel = (monroe_ionphoton_interface9_bank_bus_adr[13:9] == 4'd14);
assign monroe_ionphoton_csrbank9_pll_reset0_r = monroe_ionphoton_interface9_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank9_pll_reset0_re = ((monroe_ionphoton_csrbank9_sel & monroe_ionphoton_interface9_bank_bus_we) & (monroe_ionphoton_interface9_bank_bus_adr[0] == 1'd0));
assign monroe_ionphoton_csrbank9_pll_locked_r = monroe_ionphoton_interface9_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank9_pll_locked_re = ((monroe_ionphoton_csrbank9_sel & monroe_ionphoton_interface9_bank_bus_we) & (monroe_ionphoton_interface9_bank_bus_adr[0] == 1'd1));
assign monroe_ionphoton_rtio_crg_storage = monroe_ionphoton_rtio_crg_storage_full;
assign monroe_ionphoton_csrbank9_pll_reset0_w = monroe_ionphoton_rtio_crg_storage_full;
assign monroe_ionphoton_csrbank9_pll_locked_w = monroe_ionphoton_rtio_crg_pll_locked_status;
assign monroe_ionphoton_csrbank10_sel = (monroe_ionphoton_interface10_bank_bus_adr[13:9] == 5'd16);
assign monroe_ionphoton_csrbank10_mon_chan_sel0_r = monroe_ionphoton_interface10_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank10_mon_chan_sel0_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 1'd0));
assign monroe_ionphoton_csrbank10_mon_probe_sel0_r = monroe_ionphoton_interface10_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank10_mon_probe_sel0_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 1'd1));
assign monroe_ionphoton_mon_value_update_r = monroe_ionphoton_interface10_bank_bus_dat_w[0];
assign monroe_ionphoton_mon_value_update_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 2'd2));
assign monroe_ionphoton_csrbank10_mon_value_r = monroe_ionphoton_interface10_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank10_mon_value_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 2'd3));
assign monroe_ionphoton_csrbank10_inj_chan_sel0_r = monroe_ionphoton_interface10_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank10_inj_chan_sel0_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 3'd4));
assign monroe_ionphoton_csrbank10_inj_override_sel0_r = monroe_ionphoton_interface10_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank10_inj_override_sel0_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 3'd5));
assign monroe_ionphoton_inj_value_r = monroe_ionphoton_interface10_bank_bus_dat_w[0];
assign monroe_ionphoton_inj_value_re = ((monroe_ionphoton_csrbank10_sel & monroe_ionphoton_interface10_bank_bus_we) & (monroe_ionphoton_interface10_bank_bus_adr[2:0] == 3'd6));
assign monroe_ionphoton_mon_chan_sel_storage = monroe_ionphoton_mon_chan_sel_storage_full[5:0];
assign monroe_ionphoton_csrbank10_mon_chan_sel0_w = monroe_ionphoton_mon_chan_sel_storage_full[5:0];
assign monroe_ionphoton_mon_probe_sel_storage = monroe_ionphoton_mon_probe_sel_storage_full;
assign monroe_ionphoton_csrbank10_mon_probe_sel0_w = monroe_ionphoton_mon_probe_sel_storage_full;
assign monroe_ionphoton_csrbank10_mon_value_w = monroe_ionphoton_mon_status;
assign monroe_ionphoton_inj_chan_sel_storage = monroe_ionphoton_inj_chan_sel_storage_full[5:0];
assign monroe_ionphoton_csrbank10_inj_chan_sel0_w = monroe_ionphoton_inj_chan_sel_storage_full[5:0];
assign monroe_ionphoton_inj_override_sel_storage = monroe_ionphoton_inj_override_sel_storage_full[1:0];
assign monroe_ionphoton_csrbank10_inj_override_sel0_w = monroe_ionphoton_inj_override_sel_storage_full[1:0];
assign monroe_ionphoton_csrbank11_sel = (monroe_ionphoton_interface11_bank_bus_adr[13:9] == 4'd8);
assign monroe_ionphoton_csrbank11_bitbang0_r = monroe_ionphoton_interface11_bank_bus_dat_w[3:0];
assign monroe_ionphoton_csrbank11_bitbang0_re = ((monroe_ionphoton_csrbank11_sel & monroe_ionphoton_interface11_bank_bus_we) & (monroe_ionphoton_interface11_bank_bus_adr[1:0] == 1'd0));
assign monroe_ionphoton_csrbank11_miso_r = monroe_ionphoton_interface11_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank11_miso_re = ((monroe_ionphoton_csrbank11_sel & monroe_ionphoton_interface11_bank_bus_we) & (monroe_ionphoton_interface11_bank_bus_adr[1:0] == 1'd1));
assign monroe_ionphoton_csrbank11_bitbang_en0_r = monroe_ionphoton_interface11_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank11_bitbang_en0_re = ((monroe_ionphoton_csrbank11_sel & monroe_ionphoton_interface11_bank_bus_we) & (monroe_ionphoton_interface11_bank_bus_adr[1:0] == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage_full[3:0];
assign monroe_ionphoton_csrbank11_bitbang0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage_full[3:0];
assign monroe_ionphoton_csrbank11_miso_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_status;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage_full;
assign monroe_ionphoton_csrbank11_bitbang_en0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage_full;
assign monroe_ionphoton_csrbank12_sel = (monroe_ionphoton_interface12_bank_bus_adr[13:9] == 2'd3);
assign monroe_ionphoton_csrbank12_load7_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load7_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 1'd0));
assign monroe_ionphoton_csrbank12_load6_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load6_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 1'd1));
assign monroe_ionphoton_csrbank12_load5_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load5_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 2'd2));
assign monroe_ionphoton_csrbank12_load4_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load4_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 2'd3));
assign monroe_ionphoton_csrbank12_load3_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load3_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 3'd4));
assign monroe_ionphoton_csrbank12_load2_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load2_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 3'd5));
assign monroe_ionphoton_csrbank12_load1_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load1_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 3'd6));
assign monroe_ionphoton_csrbank12_load0_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_load0_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 3'd7));
assign monroe_ionphoton_csrbank12_reload7_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload7_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd8));
assign monroe_ionphoton_csrbank12_reload6_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload6_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd9));
assign monroe_ionphoton_csrbank12_reload5_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload5_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd10));
assign monroe_ionphoton_csrbank12_reload4_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload4_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd11));
assign monroe_ionphoton_csrbank12_reload3_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload3_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd12));
assign monroe_ionphoton_csrbank12_reload2_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload2_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd13));
assign monroe_ionphoton_csrbank12_reload1_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload1_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd14));
assign monroe_ionphoton_csrbank12_reload0_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_reload0_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 4'd15));
assign monroe_ionphoton_csrbank12_en0_r = monroe_ionphoton_interface12_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank12_en0_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd16));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_r = monroe_ionphoton_interface12_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd17));
assign monroe_ionphoton_csrbank12_value7_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value7_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd18));
assign monroe_ionphoton_csrbank12_value6_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value6_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd19));
assign monroe_ionphoton_csrbank12_value5_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value5_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd20));
assign monroe_ionphoton_csrbank12_value4_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value4_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd21));
assign monroe_ionphoton_csrbank12_value3_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value3_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd22));
assign monroe_ionphoton_csrbank12_value2_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value2_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd23));
assign monroe_ionphoton_csrbank12_value1_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value1_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd24));
assign monroe_ionphoton_csrbank12_value0_r = monroe_ionphoton_interface12_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank12_value0_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd25));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_r = monroe_ionphoton_interface12_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd26));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_r = monroe_ionphoton_interface12_bank_bus_dat_w[0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd27));
assign monroe_ionphoton_csrbank12_ev_enable0_r = monroe_ionphoton_interface12_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank12_ev_enable0_re = ((monroe_ionphoton_csrbank12_sel & monroe_ionphoton_interface12_bank_bus_we) & (monroe_ionphoton_interface12_bank_bus_adr[4:0] == 5'd28));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[63:0];
assign monroe_ionphoton_csrbank12_load7_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[63:56];
assign monroe_ionphoton_csrbank12_load6_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[55:48];
assign monroe_ionphoton_csrbank12_load5_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[47:40];
assign monroe_ionphoton_csrbank12_load4_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[39:32];
assign monroe_ionphoton_csrbank12_load3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[31:24];
assign monroe_ionphoton_csrbank12_load2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[23:16];
assign monroe_ionphoton_csrbank12_load1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[15:8];
assign monroe_ionphoton_csrbank12_load0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[63:0];
assign monroe_ionphoton_csrbank12_reload7_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[63:56];
assign monroe_ionphoton_csrbank12_reload6_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[55:48];
assign monroe_ionphoton_csrbank12_reload5_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[47:40];
assign monroe_ionphoton_csrbank12_reload4_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[39:32];
assign monroe_ionphoton_csrbank12_reload3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[31:24];
assign monroe_ionphoton_csrbank12_reload2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[23:16];
assign monroe_ionphoton_csrbank12_reload1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[15:8];
assign monroe_ionphoton_csrbank12_reload0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage_full;
assign monroe_ionphoton_csrbank12_en0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage_full;
assign monroe_ionphoton_csrbank12_value7_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[63:56];
assign monroe_ionphoton_csrbank12_value6_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[55:48];
assign monroe_ionphoton_csrbank12_value5_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[47:40];
assign monroe_ionphoton_csrbank12_value4_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[39:32];
assign monroe_ionphoton_csrbank12_value3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[31:24];
assign monroe_ionphoton_csrbank12_value2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[23:16];
assign monroe_ionphoton_csrbank12_value1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[15:8];
assign monroe_ionphoton_csrbank12_value0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage_full;
assign monroe_ionphoton_csrbank12_ev_enable0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage_full;
assign monroe_ionphoton_csrbank13_sel = (monroe_ionphoton_interface13_bank_bus_adr[13:9] == 3'd4);
assign monroe_ionphoton_csrbank13_enable_null0_r = monroe_ionphoton_interface13_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank13_enable_null0_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 1'd0));
assign monroe_ionphoton_csrbank13_enable_prog0_r = monroe_ionphoton_interface13_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank13_enable_prog0_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 1'd1));
assign monroe_ionphoton_csrbank13_prog_address3_r = monroe_ionphoton_interface13_bank_bus_dat_w[5:0];
assign monroe_ionphoton_csrbank13_prog_address3_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 2'd2));
assign monroe_ionphoton_csrbank13_prog_address2_r = monroe_ionphoton_interface13_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank13_prog_address2_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 2'd3));
assign monroe_ionphoton_csrbank13_prog_address1_r = monroe_ionphoton_interface13_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank13_prog_address1_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 3'd4));
assign monroe_ionphoton_csrbank13_prog_address0_r = monroe_ionphoton_interface13_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank13_prog_address0_re = ((monroe_ionphoton_csrbank13_sel & monroe_ionphoton_interface13_bank_bus_we) & (monroe_ionphoton_interface13_bank_bus_adr[2:0] == 3'd5));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage_full;
assign monroe_ionphoton_csrbank13_enable_null0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage_full;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage_full;
assign monroe_ionphoton_csrbank13_enable_prog0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage_full;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[29:12];
assign monroe_ionphoton_csrbank13_prog_address3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[29:24];
assign monroe_ionphoton_csrbank13_prog_address2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[23:16];
assign monroe_ionphoton_csrbank13_prog_address1_w = {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[15:12], {4{1'd0}}};
assign monroe_ionphoton_csrbank13_prog_address0_w = 1'd0;
assign monroe_ionphoton_csrbank14_sel = (monroe_ionphoton_interface14_bank_bus_adr[13:9] == 1'd1);
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_r = monroe_ionphoton_interface14_bank_bus_dat_w[7:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 1'd0));
assign monroe_ionphoton_csrbank14_txfull_r = monroe_ionphoton_interface14_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank14_txfull_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 1'd1));
assign monroe_ionphoton_csrbank14_rxempty_r = monroe_ionphoton_interface14_bank_bus_dat_w[0];
assign monroe_ionphoton_csrbank14_rxempty_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 2'd2));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_r = monroe_ionphoton_interface14_bank_bus_dat_w[1:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 2'd3));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_r = monroe_ionphoton_interface14_bank_bus_dat_w[1:0];
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 3'd4));
assign monroe_ionphoton_csrbank14_ev_enable0_r = monroe_ionphoton_interface14_bank_bus_dat_w[1:0];
assign monroe_ionphoton_csrbank14_ev_enable0_re = ((monroe_ionphoton_csrbank14_sel & monroe_ionphoton_interface14_bank_bus_we) & (monroe_ionphoton_interface14_bank_bus_adr[2:0] == 3'd5));
assign monroe_ionphoton_csrbank14_txfull_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_txfull_status;
assign monroe_ionphoton_csrbank14_rxempty_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxempty_status;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage_full[1:0];
assign monroe_ionphoton_csrbank14_ev_enable0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage_full[1:0];
assign monroe_ionphoton_csrbank15_sel = (monroe_ionphoton_interface15_bank_bus_adr[13:9] == 1'd0);
assign monroe_ionphoton_csrbank15_tuning_word3_r = monroe_ionphoton_interface15_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank15_tuning_word3_re = ((monroe_ionphoton_csrbank15_sel & monroe_ionphoton_interface15_bank_bus_we) & (monroe_ionphoton_interface15_bank_bus_adr[1:0] == 1'd0));
assign monroe_ionphoton_csrbank15_tuning_word2_r = monroe_ionphoton_interface15_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank15_tuning_word2_re = ((monroe_ionphoton_csrbank15_sel & monroe_ionphoton_interface15_bank_bus_we) & (monroe_ionphoton_interface15_bank_bus_adr[1:0] == 1'd1));
assign monroe_ionphoton_csrbank15_tuning_word1_r = monroe_ionphoton_interface15_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank15_tuning_word1_re = ((monroe_ionphoton_csrbank15_sel & monroe_ionphoton_interface15_bank_bus_we) & (monroe_ionphoton_interface15_bank_bus_adr[1:0] == 2'd2));
assign monroe_ionphoton_csrbank15_tuning_word0_r = monroe_ionphoton_interface15_bank_bus_dat_w[7:0];
assign monroe_ionphoton_csrbank15_tuning_word0_re = ((monroe_ionphoton_csrbank15_sel & monroe_ionphoton_interface15_bank_bus_we) & (monroe_ionphoton_interface15_bank_bus_adr[1:0] == 2'd3));
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[31:0];
assign monroe_ionphoton_csrbank15_tuning_word3_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[31:24];
assign monroe_ionphoton_csrbank15_tuning_word2_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[23:16];
assign monroe_ionphoton_csrbank15_tuning_word1_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[15:8];
assign monroe_ionphoton_csrbank15_tuning_word0_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[7:0];
assign monroe_ionphoton_interface0_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface1_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface2_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface3_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface4_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface5_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface6_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface7_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface8_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface9_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface10_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface11_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface12_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface13_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface14_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface15_bank_bus_adr = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr;
assign monroe_ionphoton_interface0_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface1_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface2_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface3_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface4_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface5_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface6_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface7_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface8_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface9_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface10_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface11_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface12_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface13_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface14_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface15_bank_bus_we = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we;
assign monroe_ionphoton_interface0_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface1_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface2_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface3_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface4_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface5_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface6_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface7_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface8_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface9_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface10_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface11_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface12_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface13_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface14_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_interface15_bank_bus_dat_w = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_r = (((((((((((((((monroe_ionphoton_interface0_bank_bus_dat_r | monroe_ionphoton_interface1_bank_bus_dat_r) | monroe_ionphoton_interface2_bank_bus_dat_r) | monroe_ionphoton_interface3_bank_bus_dat_r) | monroe_ionphoton_interface4_bank_bus_dat_r) | monroe_ionphoton_interface5_bank_bus_dat_r) | monroe_ionphoton_interface6_bank_bus_dat_r) | monroe_ionphoton_interface7_bank_bus_dat_r) | monroe_ionphoton_interface8_bank_bus_dat_r) | monroe_ionphoton_interface9_bank_bus_dat_r) | monroe_ionphoton_interface10_bank_bus_dat_r) | monroe_ionphoton_interface11_bank_bus_dat_r) | monroe_ionphoton_interface12_bank_bus_dat_r) | monroe_ionphoton_interface13_bank_bus_dat_r) | monroe_ionphoton_interface14_bank_bus_dat_r) | monroe_ionphoton_interface15_bank_bus_dat_r);

// synthesis translate_off
reg dummy_d_156;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed0 <= 30'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed0 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_adr;
		end
		default: begin
			comb_rhs_array_muxed0 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_156 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_157;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed1 <= 32'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed1 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_w;
		end
		default: begin
			comb_rhs_array_muxed1 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_157 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_158;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed2 <= 4'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed2 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_sel;
		end
		default: begin
			comb_rhs_array_muxed2 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_158 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_159;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed3 <= 1'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed3 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cyc;
		end
		default: begin
			comb_rhs_array_muxed3 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_159 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_160;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed4 <= 1'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed4 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_stb;
		end
		default: begin
			comb_rhs_array_muxed4 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_160 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_161;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed5 <= 1'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed5 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_we;
		end
		default: begin
			comb_rhs_array_muxed5 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_161 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_162;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed6 <= 3'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed6 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cti;
		end
		default: begin
			comb_rhs_array_muxed6 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_162 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_163;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed7 <= 2'd0;
	case (grant)
		1'd0: begin
			comb_rhs_array_muxed7 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_bte;
		end
		default: begin
			comb_rhs_array_muxed7 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_163 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_164;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed8 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record0_writable;
		end
		1'd1: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record1_writable;
		end
		2'd2: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record2_writable;
		end
		2'd3: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record3_writable;
		end
		3'd4: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record4_writable;
		end
		3'd5: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record5_writable;
		end
		3'd6: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record6_writable;
		end
		default: begin
			comb_rhs_array_muxed8 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_record7_writable;
		end
	endcase
// synthesis translate_off
	dummy_d_164 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_165;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed9 <= 2'd0;
	case (monroe_ionphoton_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow0, (monroe_ionphoton_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & (~monroe_ionphoton_rtio_core_inputs_overflow0))};
		end
		1'd1: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow1, (monroe_ionphoton_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & (~monroe_ionphoton_rtio_core_inputs_overflow1))};
		end
		2'd2: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow2, (monroe_ionphoton_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & (~monroe_ionphoton_rtio_core_inputs_overflow2))};
		end
		2'd3: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow3, (monroe_ionphoton_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & (~monroe_ionphoton_rtio_core_inputs_overflow3))};
		end
		3'd4: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd5: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd6: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd7: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd8: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd9: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd10: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd11: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd12: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd13: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd14: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd15: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd16: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow4, (monroe_ionphoton_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & (~monroe_ionphoton_rtio_core_inputs_overflow4))};
		end
		5'd17: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd18: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd19: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd20: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd21: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd22: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow5, (monroe_ionphoton_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & (~monroe_ionphoton_rtio_core_inputs_overflow5))};
		end
		5'd23: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd24: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd25: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd26: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd27: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd28: begin
			comb_rhs_array_muxed9 <= {monroe_ionphoton_rtio_core_inputs_overflow6, (monroe_ionphoton_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & (~monroe_ionphoton_rtio_core_inputs_overflow6))};
		end
		5'd29: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd30: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd31: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd32: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd33: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd34: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		6'd35: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
		default: begin
			comb_rhs_array_muxed9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_165 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_166;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed10 <= 2'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed10 <= monroe_ionphoton_rtio_cri_cmd;
		end
		default: begin
			comb_rhs_array_muxed10 <= monroe_ionphoton_dma_cri_master_cri_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_166 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_167;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed11 <= 24'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed11 <= monroe_ionphoton_rtio_cri_chan_sel;
		end
		default: begin
			comb_rhs_array_muxed11 <= monroe_ionphoton_dma_cri_master_cri_chan_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_167 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_168;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed12 <= 64'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed12 <= monroe_ionphoton_rtio_cri_o_timestamp;
		end
		default: begin
			comb_rhs_array_muxed12 <= monroe_ionphoton_dma_cri_master_cri_o_timestamp;
		end
	endcase
// synthesis translate_off
	dummy_d_168 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_169;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed13 <= 512'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed13 <= monroe_ionphoton_rtio_cri_o_data;
		end
		default: begin
			comb_rhs_array_muxed13 <= monroe_ionphoton_dma_cri_master_cri_o_data;
		end
	endcase
// synthesis translate_off
	dummy_d_169 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_170;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed14 <= 8'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed14 <= monroe_ionphoton_rtio_cri_o_address;
		end
		default: begin
			comb_rhs_array_muxed14 <= monroe_ionphoton_dma_cri_master_cri_o_address;
		end
	endcase
// synthesis translate_off
	dummy_d_170 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_171;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed15 <= 64'd0;
	case (monroe_ionphoton_cri_con_storage)
		1'd0: begin
			comb_rhs_array_muxed15 <= monroe_ionphoton_rtio_cri_i_timeout;
		end
		default: begin
			comb_rhs_array_muxed15 <= monroe_ionphoton_dma_cri_master_cri_i_timeout;
		end
	endcase
// synthesis translate_off
	dummy_d_171 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_172;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed17 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed17 <= monroe_ionphoton_inj_o_sys0;
		end
		1'd1: begin
			comb_rhs_array_muxed17 <= monroe_ionphoton_inj_o_sys1;
		end
		default: begin
			comb_rhs_array_muxed17 <= monroe_ionphoton_inj_o_sys2;
		end
	endcase
// synthesis translate_off
	dummy_d_172 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_173;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed18 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed18 <= monroe_ionphoton_inj_o_sys3;
		end
		1'd1: begin
			comb_rhs_array_muxed18 <= monroe_ionphoton_inj_o_sys4;
		end
		default: begin
			comb_rhs_array_muxed18 <= monroe_ionphoton_inj_o_sys5;
		end
	endcase
// synthesis translate_off
	dummy_d_173 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_174;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed19 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed19 <= monroe_ionphoton_inj_o_sys6;
		end
		1'd1: begin
			comb_rhs_array_muxed19 <= monroe_ionphoton_inj_o_sys7;
		end
		default: begin
			comb_rhs_array_muxed19 <= monroe_ionphoton_inj_o_sys8;
		end
	endcase
// synthesis translate_off
	dummy_d_174 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_175;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed20 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed20 <= monroe_ionphoton_inj_o_sys9;
		end
		1'd1: begin
			comb_rhs_array_muxed20 <= monroe_ionphoton_inj_o_sys10;
		end
		default: begin
			comb_rhs_array_muxed20 <= monroe_ionphoton_inj_o_sys11;
		end
	endcase
// synthesis translate_off
	dummy_d_175 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_176;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed21 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed21 <= monroe_ionphoton_inj_o_sys12;
		end
		1'd1: begin
			comb_rhs_array_muxed21 <= monroe_ionphoton_inj_o_sys13;
		end
		default: begin
			comb_rhs_array_muxed21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_176 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_177;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed22 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed22 <= monroe_ionphoton_inj_o_sys14;
		end
		1'd1: begin
			comb_rhs_array_muxed22 <= monroe_ionphoton_inj_o_sys15;
		end
		default: begin
			comb_rhs_array_muxed22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_177 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_178;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed23 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed23 <= monroe_ionphoton_inj_o_sys16;
		end
		1'd1: begin
			comb_rhs_array_muxed23 <= monroe_ionphoton_inj_o_sys17;
		end
		default: begin
			comb_rhs_array_muxed23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_178 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_179;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed24 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed24 <= monroe_ionphoton_inj_o_sys18;
		end
		1'd1: begin
			comb_rhs_array_muxed24 <= monroe_ionphoton_inj_o_sys19;
		end
		default: begin
			comb_rhs_array_muxed24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_179 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_180;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed25 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed25 <= monroe_ionphoton_inj_o_sys20;
		end
		1'd1: begin
			comb_rhs_array_muxed25 <= monroe_ionphoton_inj_o_sys21;
		end
		default: begin
			comb_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_180 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_181;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed26 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed26 <= monroe_ionphoton_inj_o_sys22;
		end
		1'd1: begin
			comb_rhs_array_muxed26 <= monroe_ionphoton_inj_o_sys23;
		end
		default: begin
			comb_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_181 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_182;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed27 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed27 <= monroe_ionphoton_inj_o_sys24;
		end
		1'd1: begin
			comb_rhs_array_muxed27 <= monroe_ionphoton_inj_o_sys25;
		end
		default: begin
			comb_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_182 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_183;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed28 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed28 <= monroe_ionphoton_inj_o_sys26;
		end
		1'd1: begin
			comb_rhs_array_muxed28 <= monroe_ionphoton_inj_o_sys27;
		end
		default: begin
			comb_rhs_array_muxed28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_183 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_184;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed29 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed29 <= monroe_ionphoton_inj_o_sys28;
		end
		1'd1: begin
			comb_rhs_array_muxed29 <= monroe_ionphoton_inj_o_sys29;
		end
		default: begin
			comb_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_184 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_185;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed30 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed30 <= monroe_ionphoton_inj_o_sys30;
		end
		1'd1: begin
			comb_rhs_array_muxed30 <= monroe_ionphoton_inj_o_sys31;
		end
		default: begin
			comb_rhs_array_muxed30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_185 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_186;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed31 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed31 <= monroe_ionphoton_inj_o_sys32;
		end
		1'd1: begin
			comb_rhs_array_muxed31 <= monroe_ionphoton_inj_o_sys33;
		end
		default: begin
			comb_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_186 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_187;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed32 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed32 <= monroe_ionphoton_inj_o_sys34;
		end
		1'd1: begin
			comb_rhs_array_muxed32 <= monroe_ionphoton_inj_o_sys35;
		end
		default: begin
			comb_rhs_array_muxed32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_187 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_188;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed33 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed33 <= 1'd0;
		end
		1'd1: begin
			comb_rhs_array_muxed33 <= 1'd0;
		end
		default: begin
			comb_rhs_array_muxed33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_188 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_189;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed34 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed34 <= monroe_ionphoton_inj_o_sys36;
		end
		1'd1: begin
			comb_rhs_array_muxed34 <= monroe_ionphoton_inj_o_sys37;
		end
		default: begin
			comb_rhs_array_muxed34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_189 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_190;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed35 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed35 <= monroe_ionphoton_inj_o_sys38;
		end
		1'd1: begin
			comb_rhs_array_muxed35 <= monroe_ionphoton_inj_o_sys39;
		end
		default: begin
			comb_rhs_array_muxed35 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_190 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_191;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed36 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed36 <= monroe_ionphoton_inj_o_sys40;
		end
		1'd1: begin
			comb_rhs_array_muxed36 <= monroe_ionphoton_inj_o_sys41;
		end
		default: begin
			comb_rhs_array_muxed36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_191 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_192;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed37 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed37 <= monroe_ionphoton_inj_o_sys42;
		end
		1'd1: begin
			comb_rhs_array_muxed37 <= monroe_ionphoton_inj_o_sys43;
		end
		default: begin
			comb_rhs_array_muxed37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_192 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_193;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed38 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed38 <= monroe_ionphoton_inj_o_sys44;
		end
		1'd1: begin
			comb_rhs_array_muxed38 <= monroe_ionphoton_inj_o_sys45;
		end
		default: begin
			comb_rhs_array_muxed38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_193 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_194;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed39 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed39 <= 1'd0;
		end
		1'd1: begin
			comb_rhs_array_muxed39 <= 1'd0;
		end
		default: begin
			comb_rhs_array_muxed39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_194 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_195;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed40 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed40 <= monroe_ionphoton_inj_o_sys46;
		end
		1'd1: begin
			comb_rhs_array_muxed40 <= monroe_ionphoton_inj_o_sys47;
		end
		default: begin
			comb_rhs_array_muxed40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_195 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_196;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed41 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed41 <= monroe_ionphoton_inj_o_sys48;
		end
		1'd1: begin
			comb_rhs_array_muxed41 <= monroe_ionphoton_inj_o_sys49;
		end
		default: begin
			comb_rhs_array_muxed41 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_196 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_197;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed42 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed42 <= monroe_ionphoton_inj_o_sys50;
		end
		1'd1: begin
			comb_rhs_array_muxed42 <= monroe_ionphoton_inj_o_sys51;
		end
		default: begin
			comb_rhs_array_muxed42 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_197 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_198;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed43 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed43 <= monroe_ionphoton_inj_o_sys52;
		end
		1'd1: begin
			comb_rhs_array_muxed43 <= monroe_ionphoton_inj_o_sys53;
		end
		default: begin
			comb_rhs_array_muxed43 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_198 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_199;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed44 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed44 <= monroe_ionphoton_inj_o_sys54;
		end
		1'd1: begin
			comb_rhs_array_muxed44 <= monroe_ionphoton_inj_o_sys55;
		end
		default: begin
			comb_rhs_array_muxed44 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_199 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_200;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed45 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed45 <= 1'd0;
		end
		1'd1: begin
			comb_rhs_array_muxed45 <= 1'd0;
		end
		default: begin
			comb_rhs_array_muxed45 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_200 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_201;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed46 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed46 <= monroe_ionphoton_inj_o_sys56;
		end
		1'd1: begin
			comb_rhs_array_muxed46 <= monroe_ionphoton_inj_o_sys57;
		end
		default: begin
			comb_rhs_array_muxed46 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_201 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_202;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed47 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed47 <= monroe_ionphoton_inj_o_sys58;
		end
		1'd1: begin
			comb_rhs_array_muxed47 <= monroe_ionphoton_inj_o_sys59;
		end
		default: begin
			comb_rhs_array_muxed47 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_202 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_203;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed48 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed48 <= monroe_ionphoton_inj_o_sys60;
		end
		1'd1: begin
			comb_rhs_array_muxed48 <= monroe_ionphoton_inj_o_sys61;
		end
		default: begin
			comb_rhs_array_muxed48 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_203 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_204;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed49 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed49 <= monroe_ionphoton_inj_o_sys62;
		end
		1'd1: begin
			comb_rhs_array_muxed49 <= monroe_ionphoton_inj_o_sys63;
		end
		default: begin
			comb_rhs_array_muxed49 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_204 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_205;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed50 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed50 <= monroe_ionphoton_inj_o_sys64;
		end
		1'd1: begin
			comb_rhs_array_muxed50 <= monroe_ionphoton_inj_o_sys65;
		end
		default: begin
			comb_rhs_array_muxed50 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_205 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_206;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed51 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed51 <= monroe_ionphoton_inj_o_sys66;
		end
		1'd1: begin
			comb_rhs_array_muxed51 <= monroe_ionphoton_inj_o_sys67;
		end
		default: begin
			comb_rhs_array_muxed51 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_206 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_207;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed52 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed52 <= monroe_ionphoton_inj_o_sys68;
		end
		1'd1: begin
			comb_rhs_array_muxed52 <= monroe_ionphoton_inj_o_sys69;
		end
		default: begin
			comb_rhs_array_muxed52 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_207 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_208;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed53 <= 1'd0;
	case (monroe_ionphoton_inj_override_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed53 <= 1'd0;
		end
		1'd1: begin
			comb_rhs_array_muxed53 <= 1'd0;
		end
		default: begin
			comb_rhs_array_muxed53 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_208 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_209;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed16 <= 1'd0;
	case (monroe_ionphoton_inj_chan_sel_storage)
		1'd0: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed17;
		end
		1'd1: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed18;
		end
		2'd2: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed19;
		end
		2'd3: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed20;
		end
		3'd4: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed21;
		end
		3'd5: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed22;
		end
		3'd6: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed23;
		end
		3'd7: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed24;
		end
		4'd8: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed25;
		end
		4'd9: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed26;
		end
		4'd10: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed27;
		end
		4'd11: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed28;
		end
		4'd12: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed29;
		end
		4'd13: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed30;
		end
		4'd14: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed31;
		end
		4'd15: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed32;
		end
		5'd16: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed33;
		end
		5'd17: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed34;
		end
		5'd18: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed35;
		end
		5'd19: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed36;
		end
		5'd20: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed37;
		end
		5'd21: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed38;
		end
		5'd22: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed39;
		end
		5'd23: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed40;
		end
		5'd24: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed41;
		end
		5'd25: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed42;
		end
		5'd26: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed43;
		end
		5'd27: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed44;
		end
		5'd28: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed45;
		end
		5'd29: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed46;
		end
		5'd30: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed47;
		end
		5'd31: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed48;
		end
		6'd32: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed49;
		end
		6'd33: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed50;
		end
		6'd34: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed51;
		end
		6'd35: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed52;
		end
		default: begin
			comb_rhs_array_muxed16 <= comb_rhs_array_muxed53;
		end
	endcase
// synthesis translate_off
	dummy_d_209 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_210;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed54 <= 30'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed54 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_adr;
		end
		default: begin
			comb_rhs_array_muxed54 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_210 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_211;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed55 <= 32'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed55 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_dat_w;
		end
		default: begin
			comb_rhs_array_muxed55 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_211 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_212;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed56 <= 4'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed56 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_sel;
		end
		default: begin
			comb_rhs_array_muxed56 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_212 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_213;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed57 <= 1'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed57 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cyc;
		end
		default: begin
			comb_rhs_array_muxed57 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_213 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_214;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed58 <= 1'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed58 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_stb;
		end
		default: begin
			comb_rhs_array_muxed58 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_214 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_215;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed59 <= 1'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed59 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_we;
		end
		default: begin
			comb_rhs_array_muxed59 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_we;
		end
	endcase
// synthesis translate_off
	dummy_d_215 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_216;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed60 <= 3'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed60 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_cti;
		end
		default: begin
			comb_rhs_array_muxed60 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_216 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_217;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed61 <= 2'd0;
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed61 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_wb_sdram_bte;
		end
		default: begin
			comb_rhs_array_muxed61 <= monroe_ionphoton_monroe_ionphoton_kernel_cpu_wb_sdram_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_217 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_218;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed62 <= 30'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed62 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_adr;
		end
		1'd1: begin
			comb_rhs_array_muxed62 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_adr;
		end
		default: begin
			comb_rhs_array_muxed62 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_218 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_219;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed63 <= 128'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed63 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_dat_w;
		end
		1'd1: begin
			comb_rhs_array_muxed63 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_dat_w;
		end
		default: begin
			comb_rhs_array_muxed63 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_219 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_220;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed64 <= 16'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed64 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_sel;
		end
		1'd1: begin
			comb_rhs_array_muxed64 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_sel;
		end
		default: begin
			comb_rhs_array_muxed64 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_220 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_221;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed65 <= 1'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed65 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cyc;
		end
		1'd1: begin
			comb_rhs_array_muxed65 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_cyc;
		end
		default: begin
			comb_rhs_array_muxed65 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_221 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_222;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed66 <= 1'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed66 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_stb;
		end
		1'd1: begin
			comb_rhs_array_muxed66 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_stb;
		end
		default: begin
			comb_rhs_array_muxed66 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_222 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_223;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed67 <= 1'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed67 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_we;
		end
		1'd1: begin
			comb_rhs_array_muxed67 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_we;
		end
		default: begin
			comb_rhs_array_muxed67 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_223 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_224;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed68 <= 3'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed68 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_cti;
		end
		1'd1: begin
			comb_rhs_array_muxed68 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_cti;
		end
		default: begin
			comb_rhs_array_muxed68 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_224 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_225;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed69 <= 2'd0;
	case (sdram_native_arbiter_grant)
		1'd0: begin
			comb_rhs_array_muxed69 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bridge_if_bus_bte;
		end
		1'd1: begin
			comb_rhs_array_muxed69 <= monroe_ionphoton_monroe_ionphoton_interface0_bus_bte;
		end
		default: begin
			comb_rhs_array_muxed69 <= monroe_ionphoton_monroe_ionphoton_interface1_bus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_225 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_226;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed70 <= 30'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed70 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_adr;
		end
		default: begin
			comb_rhs_array_muxed70 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_226 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_227;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed71 <= 32'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed71 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_w;
		end
		default: begin
			comb_rhs_array_muxed71 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_227 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_228;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed72 <= 4'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed72 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_sel;
		end
		default: begin
			comb_rhs_array_muxed72 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_228 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_229;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed73 <= 1'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed73 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cyc;
		end
		default: begin
			comb_rhs_array_muxed73 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_229 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_230;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed74 <= 1'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed74 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_stb;
		end
		default: begin
			comb_rhs_array_muxed74 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_230 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_231;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed75 <= 1'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed75 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_we;
		end
		default: begin
			comb_rhs_array_muxed75 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_we;
		end
	endcase
// synthesis translate_off
	dummy_d_231 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_232;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed76 <= 3'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed76 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cti;
		end
		default: begin
			comb_rhs_array_muxed76 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_232 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_233;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed77 <= 2'd0;
	case (monroe_ionphoton_grant)
		1'd0: begin
			comb_rhs_array_muxed77 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_bte;
		end
		default: begin
			comb_rhs_array_muxed77 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_233 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_234;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed0 <= 3'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			sync_t_rhs_array_muxed0 <= 3'd4;
		end
		2'd3: begin
			sync_t_rhs_array_muxed0 <= 2'd3;
		end
		3'd4: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			sync_t_rhs_array_muxed0 <= 2'd2;
		end
		3'd6: begin
			sync_t_rhs_array_muxed0 <= 3'd6;
		end
		3'd7: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd8: begin
			sync_t_rhs_array_muxed0 <= 3'd7;
		end
		4'd9: begin
			sync_t_rhs_array_muxed0 <= 1'd1;
		end
		4'd10: begin
			sync_t_rhs_array_muxed0 <= 3'd5;
		end
		4'd11: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd13: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd14: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_234 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_235;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed0 <= 3'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		2'd3: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		3'd4: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			sync_f_t_array_muxed0 <= 3'd5;
		end
		3'd6: begin
			sync_f_t_array_muxed0 <= 1'd1;
		end
		3'd7: begin
			sync_f_t_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		4'd9: begin
			sync_f_t_array_muxed0 <= 3'd6;
		end
		4'd10: begin
			sync_f_t_array_muxed0 <= 2'd2;
		end
		4'd11: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			sync_f_t_array_muxed0 <= 2'd3;
		end
		4'd13: begin
			sync_f_t_array_muxed0 <= 3'd4;
		end
		4'd14: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
		default: begin
			sync_f_t_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_235 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_236;
// synthesis translate_on
always @(*) begin
	sync_f_rhs_array_muxed0 <= 3'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3:0])
		1'd0: begin
			sync_f_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			sync_f_rhs_array_muxed0 <= 3'd7;
		end
		2'd2: begin
			sync_f_rhs_array_muxed0 <= 3'd4;
		end
		2'd3: begin
			sync_f_rhs_array_muxed0 <= 2'd3;
		end
		3'd4: begin
			sync_f_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			sync_f_rhs_array_muxed0 <= 2'd2;
		end
		3'd6: begin
			sync_f_rhs_array_muxed0 <= 3'd6;
		end
		3'd7: begin
			sync_f_rhs_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			sync_f_rhs_array_muxed0 <= 3'd7;
		end
		4'd9: begin
			sync_f_rhs_array_muxed0 <= 1'd1;
		end
		4'd10: begin
			sync_f_rhs_array_muxed0 <= 3'd5;
		end
		4'd11: begin
			sync_f_rhs_array_muxed0 <= 1'd0;
		end
		4'd12: begin
			sync_f_rhs_array_muxed0 <= 2'd3;
		end
		4'd13: begin
			sync_f_rhs_array_muxed0 <= 3'd4;
		end
		4'd14: begin
			sync_f_rhs_array_muxed0 <= 3'd7;
		end
		default: begin
			sync_f_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_236 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_237;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed0 <= 5'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4])
		1'd0: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		2'd3: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		3'd4: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			sync_rhs_array_muxed0 <= 5'd23;
		end
		3'd6: begin
			sync_rhs_array_muxed0 <= 4'd8;
		end
		3'd7: begin
			sync_rhs_array_muxed0 <= 3'd7;
		end
		4'd8: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		4'd9: begin
			sync_rhs_array_muxed0 <= 5'd27;
		end
		4'd10: begin
			sync_rhs_array_muxed0 <= 3'd4;
		end
		4'd11: begin
			sync_rhs_array_muxed0 <= 5'd20;
		end
		4'd12: begin
			sync_rhs_array_muxed0 <= 5'd24;
		end
		4'd13: begin
			sync_rhs_array_muxed0 <= 4'd12;
		end
		4'd14: begin
			sync_rhs_array_muxed0 <= 5'd28;
		end
		4'd15: begin
			sync_rhs_array_muxed0 <= 5'd28;
		end
		5'd16: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		5'd17: begin
			sync_rhs_array_muxed0 <= 5'd29;
		end
		5'd18: begin
			sync_rhs_array_muxed0 <= 2'd2;
		end
		5'd19: begin
			sync_rhs_array_muxed0 <= 5'd18;
		end
		5'd20: begin
			sync_rhs_array_muxed0 <= 5'd31;
		end
		5'd21: begin
			sync_rhs_array_muxed0 <= 4'd10;
		end
		5'd22: begin
			sync_rhs_array_muxed0 <= 5'd26;
		end
		5'd23: begin
			sync_rhs_array_muxed0 <= 4'd15;
		end
		5'd24: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		5'd25: begin
			sync_rhs_array_muxed0 <= 3'd6;
		end
		5'd26: begin
			sync_rhs_array_muxed0 <= 5'd22;
		end
		5'd27: begin
			sync_rhs_array_muxed0 <= 5'd16;
		end
		5'd28: begin
			sync_rhs_array_muxed0 <= 4'd14;
		end
		5'd29: begin
			sync_rhs_array_muxed0 <= 1'd1;
		end
		5'd30: begin
			sync_rhs_array_muxed0 <= 5'd30;
		end
		5'd31: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd32: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd33: begin
			sync_rhs_array_muxed0 <= 5'd30;
		end
		6'd34: begin
			sync_rhs_array_muxed0 <= 1'd1;
		end
		6'd35: begin
			sync_rhs_array_muxed0 <= 5'd17;
		end
		6'd36: begin
			sync_rhs_array_muxed0 <= 5'd16;
		end
		6'd37: begin
			sync_rhs_array_muxed0 <= 4'd9;
		end
		6'd38: begin
			sync_rhs_array_muxed0 <= 5'd25;
		end
		6'd39: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd40: begin
			sync_rhs_array_muxed0 <= 4'd15;
		end
		6'd41: begin
			sync_rhs_array_muxed0 <= 3'd5;
		end
		6'd42: begin
			sync_rhs_array_muxed0 <= 5'd21;
		end
		6'd43: begin
			sync_rhs_array_muxed0 <= 5'd31;
		end
		6'd44: begin
			sync_rhs_array_muxed0 <= 4'd13;
		end
		6'd45: begin
			sync_rhs_array_muxed0 <= 2'd2;
		end
		6'd46: begin
			sync_rhs_array_muxed0 <= 5'd29;
		end
		6'd47: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd48: begin
			sync_rhs_array_muxed0 <= 5'd28;
		end
		6'd49: begin
			sync_rhs_array_muxed0 <= 2'd3;
		end
		6'd50: begin
			sync_rhs_array_muxed0 <= 5'd19;
		end
		6'd51: begin
			sync_rhs_array_muxed0 <= 5'd24;
		end
		6'd52: begin
			sync_rhs_array_muxed0 <= 4'd11;
		end
		6'd53: begin
			sync_rhs_array_muxed0 <= 3'd4;
		end
		6'd54: begin
			sync_rhs_array_muxed0 <= 5'd27;
		end
		6'd55: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd56: begin
			sync_rhs_array_muxed0 <= 3'd7;
		end
		6'd57: begin
			sync_rhs_array_muxed0 <= 4'd8;
		end
		6'd58: begin
			sync_rhs_array_muxed0 <= 5'd23;
		end
		6'd59: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd60: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd61: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		6'd62: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
		default: begin
			sync_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_237 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_238;
// synthesis translate_on
always @(*) begin
	sync_f_rhs_array_muxed1 <= 6'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0])
		1'd0: begin
			sync_f_rhs_array_muxed1 <= 5'd24;
		end
		1'd1: begin
			sync_f_rhs_array_muxed1 <= 6'd34;
		end
		2'd2: begin
			sync_f_rhs_array_muxed1 <= 5'd18;
		end
		2'd3: begin
			sync_f_rhs_array_muxed1 <= 6'd49;
		end
		3'd4: begin
			sync_f_rhs_array_muxed1 <= 4'd10;
		end
		3'd5: begin
			sync_f_rhs_array_muxed1 <= 6'd41;
		end
		3'd6: begin
			sync_f_rhs_array_muxed1 <= 5'd25;
		end
		3'd7: begin
			sync_f_rhs_array_muxed1 <= 3'd7;
		end
		4'd8: begin
			sync_f_rhs_array_muxed1 <= 3'd6;
		end
		4'd9: begin
			sync_f_rhs_array_muxed1 <= 6'd37;
		end
		4'd10: begin
			sync_f_rhs_array_muxed1 <= 5'd21;
		end
		4'd11: begin
			sync_f_rhs_array_muxed1 <= 6'd52;
		end
		4'd12: begin
			sync_f_rhs_array_muxed1 <= 4'd13;
		end
		4'd13: begin
			sync_f_rhs_array_muxed1 <= 6'd44;
		end
		4'd14: begin
			sync_f_rhs_array_muxed1 <= 5'd28;
		end
		4'd15: begin
			sync_f_rhs_array_muxed1 <= 6'd40;
		end
		5'd16: begin
			sync_f_rhs_array_muxed1 <= 6'd36;
		end
		5'd17: begin
			sync_f_rhs_array_muxed1 <= 6'd35;
		end
		5'd18: begin
			sync_f_rhs_array_muxed1 <= 5'd19;
		end
		5'd19: begin
			sync_f_rhs_array_muxed1 <= 6'd50;
		end
		5'd20: begin
			sync_f_rhs_array_muxed1 <= 4'd11;
		end
		5'd21: begin
			sync_f_rhs_array_muxed1 <= 6'd42;
		end
		5'd22: begin
			sync_f_rhs_array_muxed1 <= 5'd26;
		end
		5'd23: begin
			sync_f_rhs_array_muxed1 <= 3'd5;
		end
		5'd24: begin
			sync_f_rhs_array_muxed1 <= 4'd12;
		end
		5'd25: begin
			sync_f_rhs_array_muxed1 <= 6'd38;
		end
		5'd26: begin
			sync_f_rhs_array_muxed1 <= 5'd22;
		end
		5'd27: begin
			sync_f_rhs_array_muxed1 <= 4'd9;
		end
		5'd28: begin
			sync_f_rhs_array_muxed1 <= 4'd14;
		end
		5'd29: begin
			sync_f_rhs_array_muxed1 <= 5'd17;
		end
		5'd30: begin
			sync_f_rhs_array_muxed1 <= 6'd33;
		end
		default: begin
			sync_f_rhs_array_muxed1 <= 5'd20;
		end
	endcase
// synthesis translate_off
	dummy_d_238 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_239;
// synthesis translate_on
always @(*) begin
	sync_f_rhs_array_muxed2 <= 1'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0])
		1'd0: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		1'd1: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		2'd2: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		2'd3: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd4: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		3'd5: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd6: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		3'd7: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd8: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		4'd9: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd10: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd11: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd12: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd13: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd14: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		4'd15: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd16: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd17: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd18: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd19: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd20: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd21: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd22: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd23: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd24: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd25: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd26: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd27: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd28: begin
			sync_f_rhs_array_muxed2 <= 1'd0;
		end
		5'd29: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		5'd30: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
		default: begin
			sync_f_rhs_array_muxed2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_239 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_240;
// synthesis translate_on
always @(*) begin
	sync_f_rhs_array_muxed3 <= 1'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0])
		1'd0: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		1'd1: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		2'd2: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		2'd3: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd4: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		3'd5: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd6: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		3'd7: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		4'd8: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		4'd9: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd10: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd11: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd12: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd13: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd14: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		4'd15: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd16: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd17: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd18: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd19: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd20: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd21: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd22: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd23: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd24: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd25: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd26: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd27: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd28: begin
			sync_f_rhs_array_muxed3 <= 1'd0;
		end
		5'd29: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		5'd30: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
		default: begin
			sync_f_rhs_array_muxed3 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_240 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_241;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed1 <= 4'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[7:5])
		1'd0: begin
			sync_rhs_array_muxed1 <= 3'd4;
		end
		1'd1: begin
			sync_rhs_array_muxed1 <= 4'd9;
		end
		2'd2: begin
			sync_rhs_array_muxed1 <= 3'd5;
		end
		2'd3: begin
			sync_rhs_array_muxed1 <= 2'd3;
		end
		3'd4: begin
			sync_rhs_array_muxed1 <= 2'd2;
		end
		3'd5: begin
			sync_rhs_array_muxed1 <= 4'd10;
		end
		3'd6: begin
			sync_rhs_array_muxed1 <= 3'd6;
		end
		default: begin
			sync_rhs_array_muxed1 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_241 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_242;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed2 <= 1'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[7:5])
		1'd0: begin
			sync_rhs_array_muxed2 <= 1'd1;
		end
		1'd1: begin
			sync_rhs_array_muxed2 <= 1'd0;
		end
		2'd2: begin
			sync_rhs_array_muxed2 <= 1'd0;
		end
		2'd3: begin
			sync_rhs_array_muxed2 <= 1'd0;
		end
		3'd4: begin
			sync_rhs_array_muxed2 <= 1'd1;
		end
		3'd5: begin
			sync_rhs_array_muxed2 <= 1'd0;
		end
		3'd6: begin
			sync_rhs_array_muxed2 <= 1'd0;
		end
		default: begin
			sync_rhs_array_muxed2 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_242 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_243;
// synthesis translate_on
always @(*) begin
	sync_f_rhs_array_muxed4 <= 1'd0;
	case (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[7:5])
		1'd0: begin
			sync_f_rhs_array_muxed4 <= 1'd1;
		end
		1'd1: begin
			sync_f_rhs_array_muxed4 <= 1'd0;
		end
		2'd2: begin
			sync_f_rhs_array_muxed4 <= 1'd0;
		end
		2'd3: begin
			sync_f_rhs_array_muxed4 <= 1'd1;
		end
		3'd4: begin
			sync_f_rhs_array_muxed4 <= 1'd1;
		end
		3'd5: begin
			sync_f_rhs_array_muxed4 <= 1'd0;
		end
		3'd6: begin
			sync_f_rhs_array_muxed4 <= 1'd0;
		end
		default: begin
			sync_f_rhs_array_muxed4 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_243 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_244;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed0 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r0)
		1'd0: begin
			sync_basiclowerer_array_muxed0 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed0 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed0 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed0 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed0 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed0 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed0 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed0 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed0 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed0 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed0 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed0 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed0 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed0 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed0 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed0 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed0 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed0 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed0 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed0 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed0 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed0 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed0 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed0 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed0 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed0 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed0 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed0 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed0 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed0 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed0 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed0 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed0 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed0 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed0 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed0 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed0 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_244 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_245;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed1 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r1)
		1'd0: begin
			sync_basiclowerer_array_muxed1 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed1 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed1 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed1 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed1 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed1 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed1 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed1 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed1 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed1 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed1 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed1 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed1 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed1 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed1 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed1 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed1 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed1 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed1 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed1 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed1 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed1 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed1 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed1 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed1 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed1 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed1 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed1 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed1 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed1 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed1 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed1 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed1 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed1 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed1 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed1 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed1 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_245 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_246;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed2 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r2)
		1'd0: begin
			sync_basiclowerer_array_muxed2 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed2 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed2 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed2 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed2 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed2 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed2 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed2 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed2 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed2 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed2 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed2 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed2 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed2 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed2 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed2 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed2 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed2 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed2 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed2 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed2 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed2 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed2 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed2 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed2 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed2 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed2 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed2 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed2 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed2 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed2 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed2 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed2 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed2 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed2 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed2 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed2 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_246 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_247;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed3 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r3)
		1'd0: begin
			sync_basiclowerer_array_muxed3 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed3 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed3 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed3 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed3 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed3 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed3 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed3 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed3 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed3 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed3 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed3 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed3 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed3 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed3 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed3 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed3 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed3 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed3 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed3 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed3 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed3 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed3 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed3 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed3 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed3 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed3 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed3 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed3 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed3 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed3 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed3 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed3 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed3 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed3 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed3 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed3 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_247 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_248;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed4 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r4)
		1'd0: begin
			sync_basiclowerer_array_muxed4 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed4 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed4 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed4 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed4 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed4 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed4 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed4 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed4 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed4 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed4 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed4 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed4 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed4 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed4 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed4 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed4 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed4 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed4 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed4 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed4 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed4 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed4 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed4 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed4 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed4 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed4 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed4 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed4 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed4 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed4 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed4 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed4 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed4 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed4 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed4 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed4 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_248 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_249;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed5 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r5)
		1'd0: begin
			sync_basiclowerer_array_muxed5 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed5 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed5 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed5 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed5 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed5 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed5 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed5 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed5 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed5 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed5 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed5 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed5 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed5 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed5 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed5 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed5 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed5 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed5 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed5 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed5 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed5 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed5 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed5 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed5 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed5 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed5 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed5 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed5 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed5 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed5 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed5 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed5 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed5 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed5 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed5 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed5 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_249 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_250;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed6 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r6)
		1'd0: begin
			sync_basiclowerer_array_muxed6 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed6 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed6 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed6 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed6 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed6 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed6 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed6 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed6 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed6 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed6 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed6 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed6 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed6 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed6 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed6 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed6 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed6 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed6 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed6 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed6 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed6 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed6 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed6 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed6 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed6 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed6 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed6 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed6 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed6 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed6 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed6 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed6 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed6 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed6 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed6 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed6 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_250 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_251;
// synthesis translate_on
always @(*) begin
	sync_basiclowerer_array_muxed7 <= 1'd0;
	case (monroe_ionphoton_rtio_core_outputs_channel_r7)
		1'd0: begin
			sync_basiclowerer_array_muxed7 <= inout_8x0_inout_8x0_ointerface0_busy;
		end
		1'd1: begin
			sync_basiclowerer_array_muxed7 <= inout_8x1_inout_8x1_ointerface1_busy;
		end
		2'd2: begin
			sync_basiclowerer_array_muxed7 <= inout_8x2_inout_8x2_ointerface2_busy;
		end
		2'd3: begin
			sync_basiclowerer_array_muxed7 <= inout_8x3_inout_8x3_ointerface3_busy;
		end
		3'd4: begin
			sync_basiclowerer_array_muxed7 <= output_8x0_busy;
		end
		3'd5: begin
			sync_basiclowerer_array_muxed7 <= output_8x1_busy;
		end
		3'd6: begin
			sync_basiclowerer_array_muxed7 <= output_8x2_busy;
		end
		3'd7: begin
			sync_basiclowerer_array_muxed7 <= output_8x3_busy;
		end
		4'd8: begin
			sync_basiclowerer_array_muxed7 <= output_8x4_busy;
		end
		4'd9: begin
			sync_basiclowerer_array_muxed7 <= output_8x5_busy;
		end
		4'd10: begin
			sync_basiclowerer_array_muxed7 <= output_8x6_busy;
		end
		4'd11: begin
			sync_basiclowerer_array_muxed7 <= output_8x7_busy;
		end
		4'd12: begin
			sync_basiclowerer_array_muxed7 <= output_8x8_busy;
		end
		4'd13: begin
			sync_basiclowerer_array_muxed7 <= output_8x9_busy;
		end
		4'd14: begin
			sync_basiclowerer_array_muxed7 <= output_8x10_busy;
		end
		4'd15: begin
			sync_basiclowerer_array_muxed7 <= output_8x11_busy;
		end
		5'd16: begin
			sync_basiclowerer_array_muxed7 <= spimaster0_ointerface0_busy;
		end
		5'd17: begin
			sync_basiclowerer_array_muxed7 <= output_8x12_busy;
		end
		5'd18: begin
			sync_basiclowerer_array_muxed7 <= output_8x13_busy;
		end
		5'd19: begin
			sync_basiclowerer_array_muxed7 <= output_8x14_busy;
		end
		5'd20: begin
			sync_basiclowerer_array_muxed7 <= output_8x15_busy;
		end
		5'd21: begin
			sync_basiclowerer_array_muxed7 <= output_8x16_busy;
		end
		5'd22: begin
			sync_basiclowerer_array_muxed7 <= spimaster1_ointerface1_busy;
		end
		5'd23: begin
			sync_basiclowerer_array_muxed7 <= output_8x17_busy;
		end
		5'd24: begin
			sync_basiclowerer_array_muxed7 <= output_8x18_busy;
		end
		5'd25: begin
			sync_basiclowerer_array_muxed7 <= output_8x19_busy;
		end
		5'd26: begin
			sync_basiclowerer_array_muxed7 <= output_8x20_busy;
		end
		5'd27: begin
			sync_basiclowerer_array_muxed7 <= output_8x21_busy;
		end
		5'd28: begin
			sync_basiclowerer_array_muxed7 <= spimaster2_ointerface2_busy;
		end
		5'd29: begin
			sync_basiclowerer_array_muxed7 <= output_8x22_busy;
		end
		5'd30: begin
			sync_basiclowerer_array_muxed7 <= output_8x23_busy;
		end
		5'd31: begin
			sync_basiclowerer_array_muxed7 <= output_8x24_busy;
		end
		6'd32: begin
			sync_basiclowerer_array_muxed7 <= output_8x25_busy;
		end
		6'd33: begin
			sync_basiclowerer_array_muxed7 <= output_8x26_busy;
		end
		6'd34: begin
			sync_basiclowerer_array_muxed7 <= output0_busy;
		end
		6'd35: begin
			sync_basiclowerer_array_muxed7 <= output1_busy;
		end
		default: begin
			sync_basiclowerer_array_muxed7 <= busy;
		end
	endcase
// synthesis translate_off
	dummy_d_251 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_252;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed1 <= 8'd0;
	case (inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed1 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed1 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed1 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed1 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed1 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed1 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed1 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed1 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_252 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_253;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed2 <= 7'd0;
	case (inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed2 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed2 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed2 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed2 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed2 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed2 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed2 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed2 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_253 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_254;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed3 <= 8'd0;
	case (inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed3 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed3 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed3 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed3 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed3 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed3 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed3 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed3 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_254 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_255;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed4 <= 7'd0;
	case (inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed4 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed4 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed4 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed4 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed4 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed4 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed4 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed4 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_255 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_256;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed5 <= 8'd0;
	case (inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed5 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed5 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed5 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed5 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed5 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed5 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed5 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed5 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_256 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_257;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed6 <= 7'd0;
	case (inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed6 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed6 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed6 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed6 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed6 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed6 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed6 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_257 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_258;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed7 <= 8'd0;
	case (inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed7 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed7 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed7 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed7 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed7 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed7 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed7 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed7 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_258 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_259;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed8 <= 7'd0;
	case (inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed8 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed8 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed8 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed8 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed8 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed8 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed8 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed8 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_259 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_260;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed9 <= 8'd0;
	case (output_8x0_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed9 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed9 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed9 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed9 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed9 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed9 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed9 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed9 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_260 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_261;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed10 <= 7'd0;
	case (output_8x0_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed10 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed10 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed10 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed10 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed10 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed10 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed10 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed10 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_261 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_262;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed11 <= 8'd0;
	case (output_8x1_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed11 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed11 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed11 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed11 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed11 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed11 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed11 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed11 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_262 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_263;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed12 <= 7'd0;
	case (output_8x1_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed12 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed12 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed12 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed12 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed12 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed12 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed12 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_263 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_264;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed13 <= 8'd0;
	case (output_8x2_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed13 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed13 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed13 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed13 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed13 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed13 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed13 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed13 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_264 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_265;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed14 <= 7'd0;
	case (output_8x2_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed14 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed14 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed14 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed14 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed14 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed14 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed14 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed14 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_265 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_266;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed15 <= 8'd0;
	case (output_8x3_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed15 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed15 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed15 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed15 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed15 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed15 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed15 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed15 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_266 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_267;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed16 <= 7'd0;
	case (output_8x3_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed16 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed16 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed16 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed16 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed16 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed16 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed16 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed16 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_267 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_268;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed17 <= 8'd0;
	case (output_8x4_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed17 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed17 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed17 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed17 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed17 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed17 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed17 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed17 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_268 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_269;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed18 <= 7'd0;
	case (output_8x4_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed18 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed18 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed18 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed18 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed18 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed18 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed18 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed18 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_269 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_270;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed19 <= 8'd0;
	case (output_8x5_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed19 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed19 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed19 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed19 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed19 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed19 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed19 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed19 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_270 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_271;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed20 <= 7'd0;
	case (output_8x5_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed20 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed20 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed20 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed20 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed20 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed20 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed20 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_271 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_272;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed21 <= 8'd0;
	case (output_8x6_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed21 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed21 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed21 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed21 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed21 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed21 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed21 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed21 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_272 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_273;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed22 <= 7'd0;
	case (output_8x6_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed22 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed22 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed22 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed22 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed22 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed22 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed22 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed22 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_273 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_274;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed23 <= 8'd0;
	case (output_8x7_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed23 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed23 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed23 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed23 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed23 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed23 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed23 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed23 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_274 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_275;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed24 <= 7'd0;
	case (output_8x7_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed24 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed24 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed24 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed24 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed24 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed24 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed24 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed24 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_275 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_276;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed25 <= 8'd0;
	case (output_8x8_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed25 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed25 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed25 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed25 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed25 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed25 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed25 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed25 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_276 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_277;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed26 <= 7'd0;
	case (output_8x8_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed26 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed26 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed26 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed26 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed26 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed26 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed26 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_277 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_278;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed27 <= 8'd0;
	case (output_8x9_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed27 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed27 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed27 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed27 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed27 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed27 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed27 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed27 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_278 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_279;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed28 <= 7'd0;
	case (output_8x9_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed28 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed28 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed28 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed28 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed28 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed28 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed28 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed28 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_279 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_280;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed29 <= 8'd0;
	case (output_8x10_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed29 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed29 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed29 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed29 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed29 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed29 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed29 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed29 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_280 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_281;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed30 <= 7'd0;
	case (output_8x10_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed30 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed30 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed30 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed30 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed30 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed30 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed30 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed30 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_281 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_282;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed31 <= 8'd0;
	case (output_8x11_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed31 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed31 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed31 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed31 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed31 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed31 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed31 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed31 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_282 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_283;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed32 <= 7'd0;
	case (output_8x11_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed32 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed32 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed32 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed32 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed32 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed32 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed32 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed32 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_283 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_284;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed33 <= 8'd0;
	case (output_8x12_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed33 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed33 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed33 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed33 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed33 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed33 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed33 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed33 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_284 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_285;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed34 <= 7'd0;
	case (output_8x12_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed34 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed34 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed34 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed34 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed34 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed34 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed34 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed34 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_285 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_286;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed35 <= 8'd0;
	case (output_8x13_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed35 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed35 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed35 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed35 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed35 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed35 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed35 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed35 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_286 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_287;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed36 <= 7'd0;
	case (output_8x13_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed36 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed36 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed36 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed36 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed36 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed36 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed36 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed36 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_287 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_288;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed37 <= 8'd0;
	case (output_8x14_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed37 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed37 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed37 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed37 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed37 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed37 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed37 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed37 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_288 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_289;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed38 <= 7'd0;
	case (output_8x14_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed38 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed38 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed38 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed38 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed38 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed38 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed38 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed38 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_289 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_290;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed39 <= 8'd0;
	case (output_8x15_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed39 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed39 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed39 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed39 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed39 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed39 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed39 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed39 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_290 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_291;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed40 <= 7'd0;
	case (output_8x15_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed40 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed40 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed40 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed40 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed40 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed40 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed40 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed40 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_291 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_292;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed41 <= 8'd0;
	case (output_8x16_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed41 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed41 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed41 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed41 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed41 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed41 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed41 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed41 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_292 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_293;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed42 <= 7'd0;
	case (output_8x16_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed42 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed42 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed42 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed42 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed42 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed42 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed42 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed42 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_293 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_294;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed43 <= 8'd0;
	case (output_8x17_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed43 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed43 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed43 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed43 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed43 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed43 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed43 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed43 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_294 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_295;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed44 <= 7'd0;
	case (output_8x17_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed44 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed44 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed44 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed44 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed44 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed44 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed44 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed44 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_295 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_296;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed45 <= 8'd0;
	case (output_8x18_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed45 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed45 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed45 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed45 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed45 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed45 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed45 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed45 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_296 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_297;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed46 <= 7'd0;
	case (output_8x18_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed46 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed46 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed46 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed46 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed46 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed46 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed46 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed46 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_297 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_298;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed47 <= 8'd0;
	case (output_8x19_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed47 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed47 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed47 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed47 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed47 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed47 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed47 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed47 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_298 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_299;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed48 <= 7'd0;
	case (output_8x19_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed48 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed48 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed48 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed48 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed48 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed48 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed48 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed48 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_299 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_300;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed49 <= 8'd0;
	case (output_8x20_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed49 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed49 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed49 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed49 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed49 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed49 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed49 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed49 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_300 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_301;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed50 <= 7'd0;
	case (output_8x20_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed50 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed50 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed50 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed50 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed50 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed50 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed50 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed50 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_301 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_302;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed51 <= 8'd0;
	case (output_8x21_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed51 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed51 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed51 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed51 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed51 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed51 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed51 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed51 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_302 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_303;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed52 <= 7'd0;
	case (output_8x21_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed52 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed52 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed52 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed52 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed52 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed52 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed52 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed52 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_303 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_304;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed53 <= 8'd0;
	case (output_8x22_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed53 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed53 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed53 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed53 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed53 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed53 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed53 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed53 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_304 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_305;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed54 <= 7'd0;
	case (output_8x22_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed54 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed54 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed54 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed54 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed54 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed54 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed54 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed54 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_305 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_306;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed55 <= 8'd0;
	case (output_8x23_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed55 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed55 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed55 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed55 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed55 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed55 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed55 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed55 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_306 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_307;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed56 <= 7'd0;
	case (output_8x23_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed56 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed56 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed56 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed56 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed56 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed56 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed56 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed56 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_307 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_308;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed57 <= 8'd0;
	case (output_8x24_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed57 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed57 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed57 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed57 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed57 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed57 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed57 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed57 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_308 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_309;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed58 <= 7'd0;
	case (output_8x24_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed58 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed58 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed58 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed58 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed58 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed58 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed58 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed58 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_309 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_310;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed59 <= 8'd0;
	case (output_8x25_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed59 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed59 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed59 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed59 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed59 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed59 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed59 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed59 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_310 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_311;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed60 <= 7'd0;
	case (output_8x25_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed60 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed60 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed60 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed60 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed60 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed60 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed60 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed60 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_311 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_312;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed61 <= 8'd0;
	case (output_8x26_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed61 <= 8'd255;
		end
		1'd1: begin
			sync_f_t_array_muxed61 <= 8'd254;
		end
		2'd2: begin
			sync_f_t_array_muxed61 <= 8'd252;
		end
		2'd3: begin
			sync_f_t_array_muxed61 <= 8'd248;
		end
		3'd4: begin
			sync_f_t_array_muxed61 <= 8'd240;
		end
		3'd5: begin
			sync_f_t_array_muxed61 <= 8'd224;
		end
		3'd6: begin
			sync_f_t_array_muxed61 <= 8'd192;
		end
		default: begin
			sync_f_t_array_muxed61 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_312 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_313;
// synthesis translate_on
always @(*) begin
	sync_f_t_array_muxed62 <= 7'd0;
	case (output_8x26_fine_ts)
		1'd0: begin
			sync_f_t_array_muxed62 <= 1'd0;
		end
		1'd1: begin
			sync_f_t_array_muxed62 <= 1'd1;
		end
		2'd2: begin
			sync_f_t_array_muxed62 <= 2'd3;
		end
		2'd3: begin
			sync_f_t_array_muxed62 <= 3'd7;
		end
		3'd4: begin
			sync_f_t_array_muxed62 <= 4'd15;
		end
		3'd5: begin
			sync_f_t_array_muxed62 <= 5'd31;
		end
		3'd6: begin
			sync_f_t_array_muxed62 <= 6'd63;
		end
		default: begin
			sync_f_t_array_muxed62 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_313 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_314;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed3 <= 61'd0;
	case (monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			sync_rhs_array_muxed3 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_314 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_315;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed4 <= 61'd0;
	case (monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_plus_one)
		1'd0: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			sync_rhs_array_muxed4 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_315 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_316;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed1 <= 32'd0;
	case (monroe_ionphoton_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record0_fifo_out_data;
		end
		1'd1: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record1_fifo_out_data;
		end
		2'd2: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record2_fifo_out_data;
		end
		2'd3: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record3_fifo_out_data;
		end
		3'd4: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd5: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd6: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd7: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd8: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd9: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd10: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd11: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd12: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd13: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd14: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd15: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd16: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record4_fifo_out_data;
		end
		5'd17: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd18: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd19: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd20: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd21: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd22: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record5_fifo_out_data;
		end
		5'd23: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd24: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd25: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd26: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd27: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd28: begin
			sync_t_rhs_array_muxed1 <= monroe_ionphoton_rtio_core_inputs_record6_fifo_out_data;
		end
		5'd29: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd30: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd31: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd32: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd33: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd34: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		6'd35: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed1 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_316 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_317;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed2 <= 65'd0;
	case (monroe_ionphoton_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			sync_t_rhs_array_muxed2 <= (monroe_ionphoton_rtio_core_inputs_record0_fifo_out_timestamp <<< 1'd0);
		end
		1'd1: begin
			sync_t_rhs_array_muxed2 <= (monroe_ionphoton_rtio_core_inputs_record1_fifo_out_timestamp <<< 1'd0);
		end
		2'd2: begin
			sync_t_rhs_array_muxed2 <= (monroe_ionphoton_rtio_core_inputs_record2_fifo_out_timestamp <<< 1'd0);
		end
		2'd3: begin
			sync_t_rhs_array_muxed2 <= (monroe_ionphoton_rtio_core_inputs_record3_fifo_out_timestamp <<< 1'd0);
		end
		3'd4: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		3'd5: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		3'd6: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		3'd7: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd8: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd9: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd10: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd11: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd12: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd13: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd14: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		4'd15: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd16: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd17: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd18: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd19: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd20: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd21: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd22: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd23: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd24: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd25: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd26: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd27: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd28: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd29: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd30: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		5'd31: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd32: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd33: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd34: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		6'd35: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed2 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_317 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_318;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed5 <= 32'd0;
	case (monroe_ionphoton_monroe_ionphoton_mailbox_i1_adr[1:0])
		1'd0: begin
			sync_rhs_array_muxed5 <= monroe_ionphoton_monroe_ionphoton_mailbox0;
		end
		1'd1: begin
			sync_rhs_array_muxed5 <= monroe_ionphoton_monroe_ionphoton_mailbox1;
		end
		default: begin
			sync_rhs_array_muxed5 <= monroe_ionphoton_monroe_ionphoton_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_318 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_319;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed6 <= 32'd0;
	case (monroe_ionphoton_monroe_ionphoton_mailbox_i2_adr[1:0])
		1'd0: begin
			sync_rhs_array_muxed6 <= monroe_ionphoton_monroe_ionphoton_mailbox0;
		end
		1'd1: begin
			sync_rhs_array_muxed6 <= monroe_ionphoton_monroe_ionphoton_mailbox1;
		end
		default: begin
			sync_rhs_array_muxed6 <= monroe_ionphoton_monroe_ionphoton_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_319 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_320;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed4 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed4 <= monroe_ionphoton_mon_bussynchronizer0_o;
		end
		default: begin
			sync_t_rhs_array_muxed4 <= monroe_ionphoton_mon_bussynchronizer1_o;
		end
	endcase
// synthesis translate_off
	dummy_d_320 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_321;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed5 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed5 <= monroe_ionphoton_mon_bussynchronizer2_o;
		end
		default: begin
			sync_t_rhs_array_muxed5 <= monroe_ionphoton_mon_bussynchronizer3_o;
		end
	endcase
// synthesis translate_off
	dummy_d_321 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_322;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed6 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed6 <= monroe_ionphoton_mon_bussynchronizer4_o;
		end
		default: begin
			sync_t_rhs_array_muxed6 <= monroe_ionphoton_mon_bussynchronizer5_o;
		end
	endcase
// synthesis translate_off
	dummy_d_322 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_323;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed7 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed7 <= monroe_ionphoton_mon_bussynchronizer6_o;
		end
		default: begin
			sync_t_rhs_array_muxed7 <= monroe_ionphoton_mon_bussynchronizer7_o;
		end
	endcase
// synthesis translate_off
	dummy_d_323 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_324;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed8 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed8 <= monroe_ionphoton_mon_bussynchronizer8_o;
		end
		default: begin
			sync_t_rhs_array_muxed8 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_324 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_325;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed9 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed9 <= monroe_ionphoton_mon_bussynchronizer9_o;
		end
		default: begin
			sync_t_rhs_array_muxed9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_325 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_326;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed10 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed10 <= monroe_ionphoton_mon_bussynchronizer10_o;
		end
		default: begin
			sync_t_rhs_array_muxed10 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_326 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_327;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed11 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed11 <= monroe_ionphoton_mon_bussynchronizer11_o;
		end
		default: begin
			sync_t_rhs_array_muxed11 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_327 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_328;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed12 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed12 <= monroe_ionphoton_mon_bussynchronizer12_o;
		end
		default: begin
			sync_t_rhs_array_muxed12 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_328 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_329;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed13 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed13 <= monroe_ionphoton_mon_bussynchronizer13_o;
		end
		default: begin
			sync_t_rhs_array_muxed13 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_329 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_330;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed14 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed14 <= monroe_ionphoton_mon_bussynchronizer14_o;
		end
		default: begin
			sync_t_rhs_array_muxed14 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_330 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_331;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed15 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed15 <= monroe_ionphoton_mon_bussynchronizer15_o;
		end
		default: begin
			sync_t_rhs_array_muxed15 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_331 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_332;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed16 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed16 <= monroe_ionphoton_mon_bussynchronizer16_o;
		end
		default: begin
			sync_t_rhs_array_muxed16 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_332 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_333;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed17 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed17 <= monroe_ionphoton_mon_bussynchronizer17_o;
		end
		default: begin
			sync_t_rhs_array_muxed17 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_333 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_334;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed18 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed18 <= monroe_ionphoton_mon_bussynchronizer18_o;
		end
		default: begin
			sync_t_rhs_array_muxed18 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_334 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_335;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed19 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed19 <= monroe_ionphoton_mon_bussynchronizer19_o;
		end
		default: begin
			sync_t_rhs_array_muxed19 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_335 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_336;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed20 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed20 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed20 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_336 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_337;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed21 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed21 <= monroe_ionphoton_mon_bussynchronizer20_o;
		end
		default: begin
			sync_t_rhs_array_muxed21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_337 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_338;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed22 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed22 <= monroe_ionphoton_mon_bussynchronizer21_o;
		end
		default: begin
			sync_t_rhs_array_muxed22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_338 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_339;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed23 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed23 <= monroe_ionphoton_mon_bussynchronizer22_o;
		end
		default: begin
			sync_t_rhs_array_muxed23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_339 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_340;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed24 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed24 <= monroe_ionphoton_mon_bussynchronizer23_o;
		end
		default: begin
			sync_t_rhs_array_muxed24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_340 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_341;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed25 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed25 <= monroe_ionphoton_mon_bussynchronizer24_o;
		end
		default: begin
			sync_t_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_341 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_342;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed26 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed26 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_342 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_343;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed27 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed27 <= monroe_ionphoton_mon_bussynchronizer25_o;
		end
		default: begin
			sync_t_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_343 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_344;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed28 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed28 <= monroe_ionphoton_mon_bussynchronizer26_o;
		end
		default: begin
			sync_t_rhs_array_muxed28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_344 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_345;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed29 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed29 <= monroe_ionphoton_mon_bussynchronizer27_o;
		end
		default: begin
			sync_t_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_345 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_346;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed30 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed30 <= monroe_ionphoton_mon_bussynchronizer28_o;
		end
		default: begin
			sync_t_rhs_array_muxed30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_346 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_347;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed31 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed31 <= monroe_ionphoton_mon_bussynchronizer29_o;
		end
		default: begin
			sync_t_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_347 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_348;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed32 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed32 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed32 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_348 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_349;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed33 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed33 <= monroe_ionphoton_mon_bussynchronizer30_o;
		end
		default: begin
			sync_t_rhs_array_muxed33 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_349 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_350;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed34 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed34 <= monroe_ionphoton_mon_bussynchronizer31_o;
		end
		default: begin
			sync_t_rhs_array_muxed34 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_350 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_351;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed35 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed35 <= monroe_ionphoton_mon_bussynchronizer32_o;
		end
		default: begin
			sync_t_rhs_array_muxed35 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_351 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_352;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed36 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed36 <= monroe_ionphoton_mon_bussynchronizer33_o;
		end
		default: begin
			sync_t_rhs_array_muxed36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_352 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_353;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed37 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed37 <= monroe_ionphoton_mon_bussynchronizer34_o;
		end
		default: begin
			sync_t_rhs_array_muxed37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_353 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_354;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed38 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed38 <= monroe_ionphoton_mon_bussynchronizer35_o;
		end
		default: begin
			sync_t_rhs_array_muxed38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_354 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_355;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed39 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed39 <= monroe_ionphoton_mon_bussynchronizer36_o;
		end
		default: begin
			sync_t_rhs_array_muxed39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_355 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_356;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed40 <= 1'd0;
	case (monroe_ionphoton_mon_probe_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed40 <= 1'd0;
		end
		default: begin
			sync_t_rhs_array_muxed40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_356 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_357;
// synthesis translate_on
always @(*) begin
	sync_t_rhs_array_muxed3 <= 1'd0;
	case (monroe_ionphoton_mon_chan_sel_storage)
		1'd0: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed4;
		end
		1'd1: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed5;
		end
		2'd2: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed6;
		end
		2'd3: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed7;
		end
		3'd4: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed8;
		end
		3'd5: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed9;
		end
		3'd6: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed10;
		end
		3'd7: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed11;
		end
		4'd8: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed12;
		end
		4'd9: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed13;
		end
		4'd10: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed14;
		end
		4'd11: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed15;
		end
		4'd12: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed16;
		end
		4'd13: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed17;
		end
		4'd14: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed18;
		end
		4'd15: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed19;
		end
		5'd16: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed20;
		end
		5'd17: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed21;
		end
		5'd18: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed22;
		end
		5'd19: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed23;
		end
		5'd20: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed24;
		end
		5'd21: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed25;
		end
		5'd22: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed26;
		end
		5'd23: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed27;
		end
		5'd24: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed28;
		end
		5'd25: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed29;
		end
		5'd26: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed30;
		end
		5'd27: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed31;
		end
		5'd28: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed32;
		end
		5'd29: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed33;
		end
		5'd30: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed34;
		end
		5'd31: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed35;
		end
		6'd32: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed36;
		end
		6'd33: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed37;
		end
		6'd34: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed38;
		end
		6'd35: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed39;
		end
		default: begin
			sync_t_rhs_array_muxed3 <= sync_t_rhs_array_muxed40;
		end
	endcase
// synthesis translate_off
	dummy_d_357 <= dummy_s;
// synthesis translate_on
end
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx = xilinxmultiregimpl0_regs1;
assign xilinxasyncresetsynchronizerimpl0 = (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_locked);
assign monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o = xilinxmultiregimpl1_regs1;
assign monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o = xilinxmultiregimpl2_regs1;
assign monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o = xilinxmultiregimpl3_regs1;
assign xilinxasyncresetsynchronizerimpl1 = (~monroe_ionphoton_monroe_ionphoton_tx_mmcm_locked);
assign xilinxasyncresetsynchronizerimpl2 = (~monroe_ionphoton_monroe_ionphoton_rx_mmcm_locked);
assign monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock1 = xilinxmultiregimpl4_regs1;
assign monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done1 = xilinxmultiregimpl5_regs1;
assign monroe_ionphoton_monroe_ionphoton_toggle_o = xilinxmultiregimpl6_regs1;
assign monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o = xilinxmultiregimpl7_regs1;
assign monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o = xilinxmultiregimpl8_regs1;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_produce_rdomain = xilinxmultiregimpl9_regs1;
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_consume_wdomain = xilinxmultiregimpl10_regs1;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_produce_rdomain = xilinxmultiregimpl11_regs1;
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_consume_wdomain = xilinxmultiregimpl12_regs1;
assign monroe_ionphoton_i2c_status1 = xilinxmultiregimpl13_regs1;
assign monroe_ionphoton_i2c_status2 = xilinxmultiregimpl14_regs1;
assign xilinxasyncresetsynchronizerimpl3 = (~monroe_ionphoton_rtio_crg_pll_locked);
assign monroe_ionphoton_rtio_crg_pll_locked_status = xilinxmultiregimpl15_regs1;
assign monroe_ionphoton_rtio_tsc_value_gray_sys = xilinxmultiregimpl16_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_produce_rdomain = xilinxmultiregimpl17_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_consume_wdomain = xilinxmultiregimpl18_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_produce_rdomain = xilinxmultiregimpl19_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_consume_wdomain = xilinxmultiregimpl20_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_produce_rdomain = xilinxmultiregimpl21_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_consume_wdomain = xilinxmultiregimpl22_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_produce_rdomain = xilinxmultiregimpl23_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_consume_wdomain = xilinxmultiregimpl24_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_produce_rdomain = xilinxmultiregimpl25_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_consume_wdomain = xilinxmultiregimpl26_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_produce_rdomain = xilinxmultiregimpl27_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_consume_wdomain = xilinxmultiregimpl28_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_produce_rdomain = xilinxmultiregimpl29_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_consume_wdomain = xilinxmultiregimpl30_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_produce_rdomain = xilinxmultiregimpl31_regs1;
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_consume_wdomain = xilinxmultiregimpl32_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_produce_rdomain = xilinxmultiregimpl33_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_consume_wdomain = xilinxmultiregimpl34_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o = xilinxmultiregimpl35_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o = xilinxmultiregimpl36_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_produce_rdomain = xilinxmultiregimpl37_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_consume_wdomain = xilinxmultiregimpl38_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o = xilinxmultiregimpl39_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o = xilinxmultiregimpl40_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_produce_rdomain = xilinxmultiregimpl41_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_consume_wdomain = xilinxmultiregimpl42_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o = xilinxmultiregimpl43_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o = xilinxmultiregimpl44_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_produce_rdomain = xilinxmultiregimpl45_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_consume_wdomain = xilinxmultiregimpl46_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o = xilinxmultiregimpl47_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o = xilinxmultiregimpl48_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_produce_rdomain = xilinxmultiregimpl49_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_consume_wdomain = xilinxmultiregimpl50_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o = xilinxmultiregimpl51_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o = xilinxmultiregimpl52_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_produce_rdomain = xilinxmultiregimpl53_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_consume_wdomain = xilinxmultiregimpl54_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o = xilinxmultiregimpl55_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o = xilinxmultiregimpl56_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_produce_rdomain = xilinxmultiregimpl57_regs1;
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_consume_wdomain = xilinxmultiregimpl58_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o = xilinxmultiregimpl59_regs1;
assign monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o = xilinxmultiregimpl60_regs1;
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o = xilinxmultiregimpl61_regs1;
assign monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o = xilinxmultiregimpl62_regs1;
assign monroe_ionphoton_rtio_core_o_collision_sync_data_o = xilinxmultiregimpl63_regs1;
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o = xilinxmultiregimpl64_regs1;
assign monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o = xilinxmultiregimpl65_regs1;
assign monroe_ionphoton_rtio_core_o_busy_sync_data_o = xilinxmultiregimpl66_regs1;
assign monroe_ionphoton_mon_bussynchronizer0_o = xilinxmultiregimpl67_regs1;
assign monroe_ionphoton_mon_bussynchronizer1_o = xilinxmultiregimpl68_regs1;
assign monroe_ionphoton_mon_bussynchronizer2_o = xilinxmultiregimpl69_regs1;
assign monroe_ionphoton_mon_bussynchronizer3_o = xilinxmultiregimpl70_regs1;
assign monroe_ionphoton_mon_bussynchronizer4_o = xilinxmultiregimpl71_regs1;
assign monroe_ionphoton_mon_bussynchronizer5_o = xilinxmultiregimpl72_regs1;
assign monroe_ionphoton_mon_bussynchronizer6_o = xilinxmultiregimpl73_regs1;
assign monroe_ionphoton_mon_bussynchronizer7_o = xilinxmultiregimpl74_regs1;
assign monroe_ionphoton_mon_bussynchronizer8_o = xilinxmultiregimpl75_regs1;
assign monroe_ionphoton_mon_bussynchronizer9_o = xilinxmultiregimpl76_regs1;
assign monroe_ionphoton_mon_bussynchronizer10_o = xilinxmultiregimpl77_regs1;
assign monroe_ionphoton_mon_bussynchronizer11_o = xilinxmultiregimpl78_regs1;
assign monroe_ionphoton_mon_bussynchronizer12_o = xilinxmultiregimpl79_regs1;
assign monroe_ionphoton_mon_bussynchronizer13_o = xilinxmultiregimpl80_regs1;
assign monroe_ionphoton_mon_bussynchronizer14_o = xilinxmultiregimpl81_regs1;
assign monroe_ionphoton_mon_bussynchronizer15_o = xilinxmultiregimpl82_regs1;
assign monroe_ionphoton_mon_bussynchronizer16_o = xilinxmultiregimpl83_regs1;
assign monroe_ionphoton_mon_bussynchronizer17_o = xilinxmultiregimpl84_regs1;
assign monroe_ionphoton_mon_bussynchronizer18_o = xilinxmultiregimpl85_regs1;
assign monroe_ionphoton_mon_bussynchronizer19_o = xilinxmultiregimpl86_regs1;
assign monroe_ionphoton_mon_bussynchronizer20_o = xilinxmultiregimpl87_regs1;
assign monroe_ionphoton_mon_bussynchronizer21_o = xilinxmultiregimpl88_regs1;
assign monroe_ionphoton_mon_bussynchronizer22_o = xilinxmultiregimpl89_regs1;
assign monroe_ionphoton_mon_bussynchronizer23_o = xilinxmultiregimpl90_regs1;
assign monroe_ionphoton_mon_bussynchronizer24_o = xilinxmultiregimpl91_regs1;
assign monroe_ionphoton_mon_bussynchronizer25_o = xilinxmultiregimpl92_regs1;
assign monroe_ionphoton_mon_bussynchronizer26_o = xilinxmultiregimpl93_regs1;
assign monroe_ionphoton_mon_bussynchronizer27_o = xilinxmultiregimpl94_regs1;
assign monroe_ionphoton_mon_bussynchronizer28_o = xilinxmultiregimpl95_regs1;
assign monroe_ionphoton_mon_bussynchronizer29_o = xilinxmultiregimpl96_regs1;
assign monroe_ionphoton_mon_bussynchronizer30_o = xilinxmultiregimpl97_regs1;
assign monroe_ionphoton_mon_bussynchronizer31_o = xilinxmultiregimpl98_regs1;
assign monroe_ionphoton_mon_bussynchronizer32_o = xilinxmultiregimpl99_regs1;
assign monroe_ionphoton_mon_bussynchronizer33_o = xilinxmultiregimpl100_regs1;
assign monroe_ionphoton_mon_bussynchronizer34_o = xilinxmultiregimpl101_regs1;
assign monroe_ionphoton_mon_bussynchronizer35_o = xilinxmultiregimpl102_regs1;
assign monroe_ionphoton_mon_bussynchronizer36_o = xilinxmultiregimpl103_regs1;
assign inout_8x0_inout_8x0_override_en = xilinxmultiregimpl104_regs1;
assign inout_8x0_inout_8x0_override_o = xilinxmultiregimpl105_regs1;
assign inout_8x0_inout_8x0_override_oe = xilinxmultiregimpl106_regs1;
assign inout_8x1_inout_8x1_override_en = xilinxmultiregimpl107_regs1;
assign inout_8x1_inout_8x1_override_o = xilinxmultiregimpl108_regs1;
assign inout_8x1_inout_8x1_override_oe = xilinxmultiregimpl109_regs1;
assign inout_8x2_inout_8x2_override_en = xilinxmultiregimpl110_regs1;
assign inout_8x2_inout_8x2_override_o = xilinxmultiregimpl111_regs1;
assign inout_8x2_inout_8x2_override_oe = xilinxmultiregimpl112_regs1;
assign inout_8x3_inout_8x3_override_en = xilinxmultiregimpl113_regs1;
assign inout_8x3_inout_8x3_override_o = xilinxmultiregimpl114_regs1;
assign inout_8x3_inout_8x3_override_oe = xilinxmultiregimpl115_regs1;
assign output_8x0_override_en = xilinxmultiregimpl116_regs1;
assign output_8x0_override_o = xilinxmultiregimpl117_regs1;
assign output_8x1_override_en = xilinxmultiregimpl118_regs1;
assign output_8x1_override_o = xilinxmultiregimpl119_regs1;
assign output_8x2_override_en = xilinxmultiregimpl120_regs1;
assign output_8x2_override_o = xilinxmultiregimpl121_regs1;
assign output_8x3_override_en = xilinxmultiregimpl122_regs1;
assign output_8x3_override_o = xilinxmultiregimpl123_regs1;
assign output_8x4_override_en = xilinxmultiregimpl124_regs1;
assign output_8x4_override_o = xilinxmultiregimpl125_regs1;
assign output_8x5_override_en = xilinxmultiregimpl126_regs1;
assign output_8x5_override_o = xilinxmultiregimpl127_regs1;
assign output_8x6_override_en = xilinxmultiregimpl128_regs1;
assign output_8x6_override_o = xilinxmultiregimpl129_regs1;
assign output_8x7_override_en = xilinxmultiregimpl130_regs1;
assign output_8x7_override_o = xilinxmultiregimpl131_regs1;
assign output_8x8_override_en = xilinxmultiregimpl132_regs1;
assign output_8x8_override_o = xilinxmultiregimpl133_regs1;
assign output_8x9_override_en = xilinxmultiregimpl134_regs1;
assign output_8x9_override_o = xilinxmultiregimpl135_regs1;
assign output_8x10_override_en = xilinxmultiregimpl136_regs1;
assign output_8x10_override_o = xilinxmultiregimpl137_regs1;
assign output_8x11_override_en = xilinxmultiregimpl138_regs1;
assign output_8x11_override_o = xilinxmultiregimpl139_regs1;
assign output_8x12_override_en = xilinxmultiregimpl140_regs1;
assign output_8x12_override_o = xilinxmultiregimpl141_regs1;
assign output_8x13_override_en = xilinxmultiregimpl142_regs1;
assign output_8x13_override_o = xilinxmultiregimpl143_regs1;
assign output_8x14_override_en = xilinxmultiregimpl144_regs1;
assign output_8x14_override_o = xilinxmultiregimpl145_regs1;
assign output_8x15_override_en = xilinxmultiregimpl146_regs1;
assign output_8x15_override_o = xilinxmultiregimpl147_regs1;
assign output_8x16_override_en = xilinxmultiregimpl148_regs1;
assign output_8x16_override_o = xilinxmultiregimpl149_regs1;
assign output_8x17_override_en = xilinxmultiregimpl150_regs1;
assign output_8x17_override_o = xilinxmultiregimpl151_regs1;
assign output_8x18_override_en = xilinxmultiregimpl152_regs1;
assign output_8x18_override_o = xilinxmultiregimpl153_regs1;
assign output_8x19_override_en = xilinxmultiregimpl154_regs1;
assign output_8x19_override_o = xilinxmultiregimpl155_regs1;
assign output_8x20_override_en = xilinxmultiregimpl156_regs1;
assign output_8x20_override_o = xilinxmultiregimpl157_regs1;
assign output_8x21_override_en = xilinxmultiregimpl158_regs1;
assign output_8x21_override_o = xilinxmultiregimpl159_regs1;
assign output_8x22_override_en = xilinxmultiregimpl160_regs1;
assign output_8x22_override_o = xilinxmultiregimpl161_regs1;
assign output_8x23_override_en = xilinxmultiregimpl162_regs1;
assign output_8x23_override_o = xilinxmultiregimpl163_regs1;
assign output_8x24_override_en = xilinxmultiregimpl164_regs1;
assign output_8x24_override_o = xilinxmultiregimpl165_regs1;
assign output_8x25_override_en = xilinxmultiregimpl166_regs1;
assign output_8x25_override_o = xilinxmultiregimpl167_regs1;
assign output_8x26_override_en = xilinxmultiregimpl168_regs1;
assign output_8x26_override_o = xilinxmultiregimpl169_regs1;
assign output0_override_en = xilinxmultiregimpl170_regs1;
assign output0_override_o = xilinxmultiregimpl171_regs1;
assign output1_override_en = xilinxmultiregimpl172_regs1;
assign output1_override_o = xilinxmultiregimpl173_regs1;

always @(posedge clk200_clk) begin
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_reset_counter != 1'd0)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_reset_counter <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_reset_counter - 1'd1);
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_reset_counter <= 4'd15;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ic_reset <= 1'd1;
	end
end

always @(posedge eth_rx_clk) begin
	monroe_ionphoton_monroe_ionphoton_pcs_rx_en_d <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en;
	monroe_ionphoton_monroe_ionphoton_pcs_source_stb <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_en;
	monroe_ionphoton_monroe_ionphoton_pcs_source_payload_data <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_rx_data;
	if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg) begin
		monroe_ionphoton_monroe_ionphoton_pcs_c_counter <= 3'd4;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_pcs_c_counter != 1'd0)) begin
			monroe_ionphoton_monroe_ionphoton_pcs_c_counter <= (monroe_ionphoton_monroe_ionphoton_pcs_c_counter - 1'd1);
		end
	end
	monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_i <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_i <= 1'd0;
	if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg) begin
		monroe_ionphoton_monroe_ionphoton_pcs_previous_config_reg <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg;
		if (((monroe_ionphoton_monroe_ionphoton_pcs_c_counter == 1'd1) & (monroe_ionphoton_monroe_ionphoton_pcs_previous_config_reg == monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg))) begin
			if (monroe_ionphoton_monroe_ionphoton_pcs_previous_config_reg[14]) begin
				monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_i <= 1'd1;
			end else begin
				monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_i <= 1'd1;
			end
		end
	end
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg <= 1'd0;
	if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_lsb) begin
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg_lsb <= monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d;
	end
	if (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_load_config_reg_msb) begin
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg <= {monroe_ionphoton_monroe_ionphoton_pcs_receivepath_d, monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg_lsb};
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] == 4'd15)) begin
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b <= sync_t_rhs_array_muxed0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] == 6'd48)) begin
			monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b <= sync_f_t_array_muxed0;
		end else begin
			if (((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3:0] == 3'd7) | (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[3:0] == 4'd8))) begin
				if (((((((monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 6'd35) & (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 5'd19)) & (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 4'd11)) & (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 6'd52)) & (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 6'd44)) & (monroe_ionphoton_monroe_ionphoton_pcs_receivepath_input_msb_first[9:4] != 5'd28))) begin
					monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k <= 1'd1;
				end
			end
			monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b <= sync_f_rhs_array_muxed0;
		end
	end
	monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code5b <= sync_rhs_array_muxed0;
	a7_1000basex_receivepath_state <= a7_1000basex_receivepath_next_state;
	if (monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_i) begin
		monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_i);
	end
	if (monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_i) begin
		monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_i);
	end
	if (monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_i) begin
		monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_i);
	end
	if ((monroe_ionphoton_monroe_ionphoton_phase_half == monroe_ionphoton_monroe_ionphoton_phase_half_rereg)) begin
		monroe_ionphoton_monroe_ionphoton_rx_data1 <= monroe_ionphoton_monroe_ionphoton_rx_data_half[19:10];
	end else begin
		monroe_ionphoton_monroe_ionphoton_rx_data1 <= monroe_ionphoton_monroe_ionphoton_rx_data_half[9:0];
	end
	monroe_ionphoton_monroe_ionphoton_phase_half <= (~monroe_ionphoton_monroe_ionphoton_phase_half);
	liteethmacpreamblechecker_state <= liteethmacpreamblechecker_next_state;
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_ce) begin
		monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg <= monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_next;
	end
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reset) begin
		monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_replace))) begin
		if ((monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce == 3'd4)) begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_do_read) begin
		if ((monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume == 3'd4)) begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_replace))) begin
		if ((~monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_do_read)) begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_do_read) begin
			monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level <= (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_fifo_reset) begin
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume <= 3'd0;
	end
	liteethmaccrc32checker_state <= liteethmaccrc32checker_next_state;
	if (monroe_ionphoton_monroe_ionphoton_ps_preamble_error_i) begin
		monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_i);
	end
	if (monroe_ionphoton_monroe_ionphoton_ps_crc_error_i) begin
		monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_i);
	end
	if (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_ack) begin
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_load_part) begin
		if (((monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux == 2'd3) | monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_eop)) begin
			monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux <= (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_stb & monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_ack)) begin
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_eop;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_stb & monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_ack)) begin
			monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop <= (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_eop | monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_load_part) begin
		case (monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux)
			1'd0: begin
				monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[39:30] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[29:20] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[19:10] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data[9:0] <= monroe_ionphoton_monroe_ionphoton_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next_binary;
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_seen_config_reg <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg <= 16'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_k <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code5b <= 5'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_code3b <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_receivepath_config_reg_lsb <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_source_stb <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_source_payload_data <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_rx_en_d <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_i <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_i <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_c_counter <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_previous_config_reg <= 16'd0;
		monroe_ionphoton_monroe_ionphoton_rx_data1 <= 10'd0;
		monroe_ionphoton_monroe_ionphoton_phase_half <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_crc_reg <= 32'd4294967295;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_level <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_produce <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_consume <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_eop <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_source_payload_data <= 40'd0;
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_demux <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_rx_converter_converter_strobe_all <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q_binary <= 7'd0;
		a7_1000basex_receivepath_state <= 3'd0;
		liteethmacpreamblechecker_state <= 1'd0;
		liteethmaccrc32checker_state <= 2'd0;
	end
	xilinxmultiregimpl12_regs0 <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q;
	xilinxmultiregimpl12_regs1 <= xilinxmultiregimpl12_regs0;
end

always @(posedge eth_rx_half_clk) begin
	monroe_ionphoton_monroe_ionphoton_phase_half_rereg <= monroe_ionphoton_monroe_ionphoton_phase_half;
end

always @(posedge eth_tx_clk) begin
	monroe_ionphoton_monroe_ionphoton_pcs_checker_tick <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_pcs_checker_counter == 1'd0)) begin
		monroe_ionphoton_monroe_ionphoton_pcs_checker_tick <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_pcs_checker_counter <= 20'd750000;
	end else begin
		monroe_ionphoton_monroe_ionphoton_pcs_checker_counter <= (monroe_ionphoton_monroe_ionphoton_pcs_checker_counter - 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_o) begin
		monroe_ionphoton_monroe_ionphoton_pcs_checker_ok <= 1'd1;
	end
	if (monroe_ionphoton_monroe_ionphoton_pcs_checker_tick) begin
		monroe_ionphoton_monroe_ionphoton_pcs_checker_ok <= 1'd0;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_parity <= (~monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_parity);
	if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_load_config_reg_buffer) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg_buffer <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_in <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output0 <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output1;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disparity <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_out;
	if ((monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k1 & (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 5'd28))) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b <= 6'd48;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_unbalanced <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_flip <= 1'd1;
	end else begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b <= sync_f_rhs_array_muxed1;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_unbalanced <= sync_f_rhs_array_muxed2;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_flip <= sync_f_rhs_array_muxed3;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b <= sync_rhs_array_muxed1;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_unbalanced <= sync_rhs_array_muxed2;
	if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k1) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_flip <= 1'd1;
	end else begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_flip <= sync_f_rhs_array_muxed4;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0 <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1 <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[7:5] == 3'd7)) begin
		if ((((monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 5'd17) | (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 5'd18)) | (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 5'd20))) begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0 <= 1'd1;
		end
		if ((((monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 4'd11) | (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 4'd13)) | (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_d1[4:0] == 4'd14))) begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1 <= 1'd1;
		end
		if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_k1) begin
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0 <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1 <= 1'd1;
		end
	end
	a7_1000basex_transmitpath_state <= a7_1000basex_transmitpath_next_state;
	if (monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value_ce) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type <= monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type_pcs_next_value;
	end
	monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_o;
	monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_o;
	monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_o;
	if (monroe_ionphoton_monroe_ionphoton_pcs_wait) begin
		if ((~monroe_ionphoton_monroe_ionphoton_pcs_done)) begin
			monroe_ionphoton_monroe_ionphoton_pcs_count <= (monroe_ionphoton_monroe_ionphoton_pcs_count - 1'd1);
		end
	end else begin
		monroe_ionphoton_monroe_ionphoton_pcs_count <= 21'd1250000;
	end
	a7_1000basex_fsm_state <= a7_1000basex_fsm_next_state;
	if (monroe_ionphoton_monroe_ionphoton_i) begin
		monroe_ionphoton_monroe_ionphoton_toggle_i <= (~monroe_ionphoton_monroe_ionphoton_toggle_i);
	end
	monroe_ionphoton_monroe_ionphoton_buf <= {monroe_ionphoton_monroe_ionphoton_tx_data1, monroe_ionphoton_monroe_ionphoton_buf[19:10]};
	if (monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_reset) begin
		monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter_ce) begin
			monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter <= (monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter + 1'd1);
		end
	end
	liteethmacgap_state <= liteethmacgap_next_state;
	if (monroe_ionphoton_monroe_ionphoton_preamble_inserter_clr_cnt) begin
		monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_preamble_inserter_inc_cnt) begin
			monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt <= (monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt + 1'd1);
		end
	end
	liteethmacpreambleinserter_state <= liteethmacpreambleinserter_next_state;
	if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing0) begin
		monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_crc32_inserter_is_ongoing1 & (~monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt_done))) begin
			monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt <= (monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt - monroe_ionphoton_monroe_ionphoton_crc32_inserter_source_ack);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_ce) begin
		monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg <= monroe_ionphoton_monroe_ionphoton_crc32_inserter_next;
	end
	if (monroe_ionphoton_monroe_ionphoton_crc32_inserter_reset) begin
		monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg <= 32'd4294967295;
	end
	liteethmaccrc32inserter_state <= liteethmaccrc32inserter_next_state;
	if (monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_reset) begin
		monroe_ionphoton_monroe_ionphoton_padding_inserter_counter <= 1'd0;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_padding_inserter_counter_ce) begin
			monroe_ionphoton_monroe_ionphoton_padding_inserter_counter <= (monroe_ionphoton_monroe_ionphoton_padding_inserter_counter + 1'd1);
		end
	end
	liteethmacpaddinginserter_state <= liteethmacpaddinginserter_next_state;
	if ((monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_stb & monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_ack)) begin
		if (monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_eop) begin
			monroe_ionphoton_monroe_ionphoton_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (monroe_ionphoton_monroe_ionphoton_tx_last_be_sink_payload_last_be) begin
				monroe_ionphoton_monroe_ionphoton_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_stb & monroe_ionphoton_monroe_ionphoton_tx_converter_converter_source_ack)) begin
		if (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_last) begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux <= 1'd0;
		end else begin
			monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux <= (monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux + 1'd1);
		end
	end
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_binary <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next_binary;
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_output0 <= 10'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disparity <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_disp_in <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_unbalanced <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code6b_flip <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_unbalanced <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_code4b_flip <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_alt7_rd1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_parity <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_c_type <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_transmitpath_config_reg_buffer <= 16'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_checker_counter <= 20'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_checker_tick <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_checker_ok <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_pcs_count <= 21'd1250000;
		monroe_ionphoton_monroe_ionphoton_buf <= 20'd0;
		monroe_ionphoton_monroe_ionphoton_tx_gap_inserter_counter <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_preamble_inserter_cnt <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_crc32_inserter_reg <= 32'd4294967295;
		monroe_ionphoton_monroe_ionphoton_crc32_inserter_cnt <= 2'd3;
		monroe_ionphoton_monroe_ionphoton_padding_inserter_counter <= 16'd1;
		monroe_ionphoton_monroe_ionphoton_tx_last_be_ongoing <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_tx_converter_converter_mux <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q_binary <= 7'd0;
		a7_1000basex_transmitpath_state <= 3'd0;
		a7_1000basex_fsm_state <= 2'd0;
		liteethmacgap_state <= 1'd0;
		liteethmacpreambleinserter_state <= 2'd0;
		liteethmaccrc32inserter_state <= 2'd0;
		liteethmacpaddinginserter_state <= 1'd0;
	end
	xilinxmultiregimpl1_regs0 <= monroe_ionphoton_monroe_ionphoton_pcs_seen_valid_ci_toggle_i;
	xilinxmultiregimpl1_regs1 <= xilinxmultiregimpl1_regs0;
	xilinxmultiregimpl2_regs0 <= monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_toggle_i;
	xilinxmultiregimpl2_regs1 <= xilinxmultiregimpl2_regs0;
	xilinxmultiregimpl3_regs0 <= monroe_ionphoton_monroe_ionphoton_pcs_rx_config_reg_ack_toggle_i;
	xilinxmultiregimpl3_regs1 <= xilinxmultiregimpl3_regs0;
	xilinxmultiregimpl9_regs0 <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q;
	xilinxmultiregimpl9_regs1 <= xilinxmultiregimpl9_regs0;
end

always @(posedge eth_tx_half_clk) begin
	monroe_ionphoton_monroe_ionphoton_tx_data_half <= monroe_ionphoton_monroe_ionphoton_buf;
end

always @(posedge rio_clk) begin
	inout_8x0_inout_8x0_sample <= 1'd0;
	if ((inout_8x0_inout_8x0_ointerface0_stb & inout_8x0_inout_8x0_ointerface0_address[1])) begin
		inout_8x0_inout_8x0_sensitivity <= inout_8x0_inout_8x0_ointerface0_data;
		if (inout_8x0_inout_8x0_ointerface0_address[0]) begin
			inout_8x0_inout_8x0_sample <= 1'd1;
		end
	end
	inout_8x1_inout_8x1_sample <= 1'd0;
	if ((inout_8x1_inout_8x1_ointerface1_stb & inout_8x1_inout_8x1_ointerface1_address[1])) begin
		inout_8x1_inout_8x1_sensitivity <= inout_8x1_inout_8x1_ointerface1_data;
		if (inout_8x1_inout_8x1_ointerface1_address[0]) begin
			inout_8x1_inout_8x1_sample <= 1'd1;
		end
	end
	inout_8x2_inout_8x2_sample <= 1'd0;
	if ((inout_8x2_inout_8x2_ointerface2_stb & inout_8x2_inout_8x2_ointerface2_address[1])) begin
		inout_8x2_inout_8x2_sensitivity <= inout_8x2_inout_8x2_ointerface2_data;
		if (inout_8x2_inout_8x2_ointerface2_address[0]) begin
			inout_8x2_inout_8x2_sample <= 1'd1;
		end
	end
	inout_8x3_inout_8x3_sample <= 1'd0;
	if ((inout_8x3_inout_8x3_ointerface3_stb & inout_8x3_inout_8x3_ointerface3_address[1])) begin
		inout_8x3_inout_8x3_sensitivity <= inout_8x3_inout_8x3_ointerface3_data;
		if (inout_8x3_inout_8x3_ointerface3_address[0]) begin
			inout_8x3_inout_8x3_sample <= 1'd1;
		end
	end
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
	if ((monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_re | (~monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable))) begin
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_dout <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
	monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record0_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record0_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record0_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record0_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record0_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record0_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record0_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record0_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record0_re & monroe_ionphoton_rtio_core_outputs_gates_record0_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record1_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record1_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record1_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record1_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record1_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record1_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record1_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record1_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record1_re & monroe_ionphoton_rtio_core_outputs_gates_record1_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record2_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record2_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record2_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record2_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record2_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record2_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record2_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record2_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record2_re & monroe_ionphoton_rtio_core_outputs_gates_record2_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record3_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record3_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record3_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record3_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record3_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record3_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record3_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record3_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record3_re & monroe_ionphoton_rtio_core_outputs_gates_record3_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record4_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record4_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record4_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record4_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record4_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record4_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record4_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record4_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record4_re & monroe_ionphoton_rtio_core_outputs_gates_record4_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record5_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record5_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record5_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record5_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record5_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record5_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record5_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record5_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record5_re & monroe_ionphoton_rtio_core_outputs_gates_record5_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record6_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record6_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record6_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record6_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record6_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record6_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record6_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record6_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record6_re & monroe_ionphoton_rtio_core_outputs_gates_record6_readable);
	monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel1 <= monroe_ionphoton_rtio_core_outputs_gates_record7_payload_channel0;
	monroe_ionphoton_rtio_core_outputs_gates_record7_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_gates_record7_payload_timestamp[2:0];
	monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address1 <= monroe_ionphoton_rtio_core_outputs_gates_record7_payload_address0;
	monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data1 <= monroe_ionphoton_rtio_core_outputs_gates_record7_payload_data0;
	monroe_ionphoton_rtio_core_outputs_gates_record7_seqn1 <= monroe_ionphoton_rtio_core_outputs_gates_record7_seqn0;
	monroe_ionphoton_rtio_core_outputs_gates_record7_valid <= (monroe_ionphoton_rtio_core_outputs_gates_record7_re & monroe_ionphoton_rtio_core_outputs_gates_record7_readable);
	monroe_ionphoton_rtio_core_outputs_record0_valid1 <= monroe_ionphoton_rtio_core_outputs_record40_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record0_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record40_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record40_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record0_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record40_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record0_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record40_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r0 <= monroe_ionphoton_rtio_core_outputs_record40_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r0 <= monroe_ionphoton_rtio_core_outputs_record40_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record1_valid1 <= monroe_ionphoton_rtio_core_outputs_record41_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record1_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record1_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record1_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r1 <= monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r1 <= monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record2_valid1 <= monroe_ionphoton_rtio_core_outputs_record42_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record2_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record2_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record2_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r2 <= monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r2 <= monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record3_valid1 <= monroe_ionphoton_rtio_core_outputs_record43_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record3_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record3_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record3_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r3 <= monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r3 <= monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record4_valid1 <= monroe_ionphoton_rtio_core_outputs_record44_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record4_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record4_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record4_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r4 <= monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r4 <= monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record5_valid1 <= monroe_ionphoton_rtio_core_outputs_record45_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record5_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record5_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record5_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r5 <= monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r5 <= monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record6_valid1 <= monroe_ionphoton_rtio_core_outputs_record46_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record6_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record6_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record6_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r6 <= monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r6 <= monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record7_valid1 <= monroe_ionphoton_rtio_core_outputs_record47_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record7_payload_channel3 <= monroe_ionphoton_rtio_core_outputs_record47_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1 <= monroe_ionphoton_rtio_core_outputs_record47_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record7_payload_address3 <= monroe_ionphoton_rtio_core_outputs_record47_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record7_payload_data3 <= monroe_ionphoton_rtio_core_outputs_record47_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_replace_occured_r7 <= monroe_ionphoton_rtio_core_outputs_record47_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r7 <= monroe_ionphoton_rtio_core_outputs_record47_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_collision <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_collision_channel <= 1'd0;
	if ((monroe_ionphoton_rtio_core_outputs_record0_valid1 & monroe_ionphoton_rtio_core_outputs_record0_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record1_valid1 & monroe_ionphoton_rtio_core_outputs_record1_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record2_valid1 & monroe_ionphoton_rtio_core_outputs_record2_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record3_valid1 & monroe_ionphoton_rtio_core_outputs_record3_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record4_valid1 & monroe_ionphoton_rtio_core_outputs_record4_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record5_valid1 & monroe_ionphoton_rtio_core_outputs_record5_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record6_valid1 & monroe_ionphoton_rtio_core_outputs_record6_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel3;
	end
	if ((monroe_ionphoton_rtio_core_outputs_record7_valid1 & monroe_ionphoton_rtio_core_outputs_record7_collision)) begin
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_collision_channel <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel3;
	end
	inout_8x0_inout_8x0_ointerface0_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected0 | monroe_ionphoton_rtio_core_outputs_selected1) | monroe_ionphoton_rtio_core_outputs_selected2) | monroe_ionphoton_rtio_core_outputs_selected3) | monroe_ionphoton_rtio_core_outputs_selected4) | monroe_ionphoton_rtio_core_outputs_selected5) | monroe_ionphoton_rtio_core_outputs_selected6) | monroe_ionphoton_rtio_core_outputs_selected7);
	inout_8x0_inout_8x0_ointerface0_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected0 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected1 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected2 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected3 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected4 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected5 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected6 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected7 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	inout_8x0_inout_8x0_ointerface0_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected0 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected1 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected2 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected3 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected4 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected5 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected6 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected7 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	inout_8x0_inout_8x0_ointerface0_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected0 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected1 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected2 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected3 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected4 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected5 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected6 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected7 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	inout_8x1_inout_8x1_ointerface1_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected8 | monroe_ionphoton_rtio_core_outputs_selected9) | monroe_ionphoton_rtio_core_outputs_selected10) | monroe_ionphoton_rtio_core_outputs_selected11) | monroe_ionphoton_rtio_core_outputs_selected12) | monroe_ionphoton_rtio_core_outputs_selected13) | monroe_ionphoton_rtio_core_outputs_selected14) | monroe_ionphoton_rtio_core_outputs_selected15);
	inout_8x1_inout_8x1_ointerface1_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected8 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected9 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected10 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected11 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected12 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected13 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected14 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected15 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	inout_8x1_inout_8x1_ointerface1_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected8 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected9 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected10 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected11 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected12 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected13 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected14 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected15 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	inout_8x1_inout_8x1_ointerface1_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected8 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected9 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected10 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected11 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected12 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected13 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected14 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected15 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	inout_8x2_inout_8x2_ointerface2_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected16 | monroe_ionphoton_rtio_core_outputs_selected17) | monroe_ionphoton_rtio_core_outputs_selected18) | monroe_ionphoton_rtio_core_outputs_selected19) | monroe_ionphoton_rtio_core_outputs_selected20) | monroe_ionphoton_rtio_core_outputs_selected21) | monroe_ionphoton_rtio_core_outputs_selected22) | monroe_ionphoton_rtio_core_outputs_selected23);
	inout_8x2_inout_8x2_ointerface2_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected16 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected17 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected18 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected19 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected20 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected21 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected22 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected23 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	inout_8x2_inout_8x2_ointerface2_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected16 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected17 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected18 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected19 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected20 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected21 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected22 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected23 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	inout_8x2_inout_8x2_ointerface2_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected16 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected17 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected18 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected19 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected20 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected21 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected22 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected23 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	inout_8x3_inout_8x3_ointerface3_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected24 | monroe_ionphoton_rtio_core_outputs_selected25) | monroe_ionphoton_rtio_core_outputs_selected26) | monroe_ionphoton_rtio_core_outputs_selected27) | monroe_ionphoton_rtio_core_outputs_selected28) | monroe_ionphoton_rtio_core_outputs_selected29) | monroe_ionphoton_rtio_core_outputs_selected30) | monroe_ionphoton_rtio_core_outputs_selected31);
	inout_8x3_inout_8x3_ointerface3_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected24 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected25 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected26 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected27 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected28 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected29 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected30 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected31 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	inout_8x3_inout_8x3_ointerface3_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected24 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected25 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected26 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected27 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected28 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected29 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected30 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected31 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	inout_8x3_inout_8x3_ointerface3_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected24 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected25 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected26 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected27 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected28 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected29 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected30 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected31 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x0_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected32 | monroe_ionphoton_rtio_core_outputs_selected33) | monroe_ionphoton_rtio_core_outputs_selected34) | monroe_ionphoton_rtio_core_outputs_selected35) | monroe_ionphoton_rtio_core_outputs_selected36) | monroe_ionphoton_rtio_core_outputs_selected37) | monroe_ionphoton_rtio_core_outputs_selected38) | monroe_ionphoton_rtio_core_outputs_selected39);
	output_8x0_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected32 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected33 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected34 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected35 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected36 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected37 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected38 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected39 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x0_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected32 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected33 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected34 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected35 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected36 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected37 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected38 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected39 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x1_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected40 | monroe_ionphoton_rtio_core_outputs_selected41) | monroe_ionphoton_rtio_core_outputs_selected42) | monroe_ionphoton_rtio_core_outputs_selected43) | monroe_ionphoton_rtio_core_outputs_selected44) | monroe_ionphoton_rtio_core_outputs_selected45) | monroe_ionphoton_rtio_core_outputs_selected46) | monroe_ionphoton_rtio_core_outputs_selected47);
	output_8x1_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected40 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected41 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected42 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected43 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected44 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected45 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected46 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected47 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x1_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected40 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected41 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected42 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected43 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected44 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected45 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected46 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected47 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x2_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected48 | monroe_ionphoton_rtio_core_outputs_selected49) | monroe_ionphoton_rtio_core_outputs_selected50) | monroe_ionphoton_rtio_core_outputs_selected51) | monroe_ionphoton_rtio_core_outputs_selected52) | monroe_ionphoton_rtio_core_outputs_selected53) | monroe_ionphoton_rtio_core_outputs_selected54) | monroe_ionphoton_rtio_core_outputs_selected55);
	output_8x2_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected48 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected49 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected50 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected51 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected52 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected53 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected54 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected55 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x2_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected48 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected49 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected50 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected51 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected52 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected53 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected54 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected55 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x3_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected56 | monroe_ionphoton_rtio_core_outputs_selected57) | monroe_ionphoton_rtio_core_outputs_selected58) | monroe_ionphoton_rtio_core_outputs_selected59) | monroe_ionphoton_rtio_core_outputs_selected60) | monroe_ionphoton_rtio_core_outputs_selected61) | monroe_ionphoton_rtio_core_outputs_selected62) | monroe_ionphoton_rtio_core_outputs_selected63);
	output_8x3_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected56 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected57 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected58 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected59 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected60 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected61 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected62 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected63 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x3_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected56 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected57 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected58 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected59 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected60 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected61 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected62 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected63 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x4_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected64 | monroe_ionphoton_rtio_core_outputs_selected65) | monroe_ionphoton_rtio_core_outputs_selected66) | monroe_ionphoton_rtio_core_outputs_selected67) | monroe_ionphoton_rtio_core_outputs_selected68) | monroe_ionphoton_rtio_core_outputs_selected69) | monroe_ionphoton_rtio_core_outputs_selected70) | monroe_ionphoton_rtio_core_outputs_selected71);
	output_8x4_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected64 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected65 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected66 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected67 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected68 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected69 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected70 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected71 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x4_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected64 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected65 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected66 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected67 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected68 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected69 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected70 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected71 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x5_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected72 | monroe_ionphoton_rtio_core_outputs_selected73) | monroe_ionphoton_rtio_core_outputs_selected74) | monroe_ionphoton_rtio_core_outputs_selected75) | monroe_ionphoton_rtio_core_outputs_selected76) | monroe_ionphoton_rtio_core_outputs_selected77) | monroe_ionphoton_rtio_core_outputs_selected78) | monroe_ionphoton_rtio_core_outputs_selected79);
	output_8x5_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected72 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected73 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected74 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected75 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected76 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected77 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected78 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected79 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x5_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected72 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected73 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected74 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected75 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected76 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected77 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected78 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected79 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x6_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected80 | monroe_ionphoton_rtio_core_outputs_selected81) | monroe_ionphoton_rtio_core_outputs_selected82) | monroe_ionphoton_rtio_core_outputs_selected83) | monroe_ionphoton_rtio_core_outputs_selected84) | monroe_ionphoton_rtio_core_outputs_selected85) | monroe_ionphoton_rtio_core_outputs_selected86) | monroe_ionphoton_rtio_core_outputs_selected87);
	output_8x6_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected80 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected81 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected82 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected83 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected84 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected85 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected86 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected87 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x6_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected80 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected81 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected82 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected83 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected84 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected85 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected86 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected87 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x7_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected88 | monroe_ionphoton_rtio_core_outputs_selected89) | monroe_ionphoton_rtio_core_outputs_selected90) | monroe_ionphoton_rtio_core_outputs_selected91) | monroe_ionphoton_rtio_core_outputs_selected92) | monroe_ionphoton_rtio_core_outputs_selected93) | monroe_ionphoton_rtio_core_outputs_selected94) | monroe_ionphoton_rtio_core_outputs_selected95);
	output_8x7_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected88 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected89 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected90 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected91 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected92 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected93 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected94 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected95 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x7_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected88 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected89 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected90 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected91 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected92 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected93 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected94 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected95 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x8_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected96 | monroe_ionphoton_rtio_core_outputs_selected97) | monroe_ionphoton_rtio_core_outputs_selected98) | monroe_ionphoton_rtio_core_outputs_selected99) | monroe_ionphoton_rtio_core_outputs_selected100) | monroe_ionphoton_rtio_core_outputs_selected101) | monroe_ionphoton_rtio_core_outputs_selected102) | monroe_ionphoton_rtio_core_outputs_selected103);
	output_8x8_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected96 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected97 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected98 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected99 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected100 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected101 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected102 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected103 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x8_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected96 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected97 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected98 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected99 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected100 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected101 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected102 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected103 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x9_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected104 | monroe_ionphoton_rtio_core_outputs_selected105) | monroe_ionphoton_rtio_core_outputs_selected106) | monroe_ionphoton_rtio_core_outputs_selected107) | monroe_ionphoton_rtio_core_outputs_selected108) | monroe_ionphoton_rtio_core_outputs_selected109) | monroe_ionphoton_rtio_core_outputs_selected110) | monroe_ionphoton_rtio_core_outputs_selected111);
	output_8x9_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected104 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected105 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected106 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected107 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected108 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected109 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected110 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected111 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x9_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected104 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected105 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected106 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected107 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected108 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected109 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected110 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected111 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x10_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected112 | monroe_ionphoton_rtio_core_outputs_selected113) | monroe_ionphoton_rtio_core_outputs_selected114) | monroe_ionphoton_rtio_core_outputs_selected115) | monroe_ionphoton_rtio_core_outputs_selected116) | monroe_ionphoton_rtio_core_outputs_selected117) | monroe_ionphoton_rtio_core_outputs_selected118) | monroe_ionphoton_rtio_core_outputs_selected119);
	output_8x10_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected112 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected113 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected114 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected115 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected116 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected117 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected118 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected119 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x10_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected112 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected113 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected114 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected115 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected116 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected117 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected118 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected119 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x11_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected120 | monroe_ionphoton_rtio_core_outputs_selected121) | monroe_ionphoton_rtio_core_outputs_selected122) | monroe_ionphoton_rtio_core_outputs_selected123) | monroe_ionphoton_rtio_core_outputs_selected124) | monroe_ionphoton_rtio_core_outputs_selected125) | monroe_ionphoton_rtio_core_outputs_selected126) | monroe_ionphoton_rtio_core_outputs_selected127);
	output_8x11_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected120 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected121 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected122 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected123 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected124 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected125 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected126 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected127 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x11_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected120 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected121 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected122 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected123 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected124 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected125 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected126 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected127 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	spimaster0_ointerface0_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected128 | monroe_ionphoton_rtio_core_outputs_selected129) | monroe_ionphoton_rtio_core_outputs_selected130) | monroe_ionphoton_rtio_core_outputs_selected131) | monroe_ionphoton_rtio_core_outputs_selected132) | monroe_ionphoton_rtio_core_outputs_selected133) | monroe_ionphoton_rtio_core_outputs_selected134) | monroe_ionphoton_rtio_core_outputs_selected135);
	spimaster0_ointerface0_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected128 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected129 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected130 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected131 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected132 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected133 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected134 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected135 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	spimaster0_ointerface0_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected128 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected129 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected130 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected131 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected132 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected133 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected134 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected135 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x12_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected136 | monroe_ionphoton_rtio_core_outputs_selected137) | monroe_ionphoton_rtio_core_outputs_selected138) | monroe_ionphoton_rtio_core_outputs_selected139) | monroe_ionphoton_rtio_core_outputs_selected140) | monroe_ionphoton_rtio_core_outputs_selected141) | monroe_ionphoton_rtio_core_outputs_selected142) | monroe_ionphoton_rtio_core_outputs_selected143);
	output_8x12_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected136 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected137 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected138 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected139 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected140 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected141 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected142 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected143 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x12_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected136 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected137 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected138 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected139 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected140 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected141 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected142 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected143 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x13_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected144 | monroe_ionphoton_rtio_core_outputs_selected145) | monroe_ionphoton_rtio_core_outputs_selected146) | monroe_ionphoton_rtio_core_outputs_selected147) | monroe_ionphoton_rtio_core_outputs_selected148) | monroe_ionphoton_rtio_core_outputs_selected149) | monroe_ionphoton_rtio_core_outputs_selected150) | monroe_ionphoton_rtio_core_outputs_selected151);
	output_8x13_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected144 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected145 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected146 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected147 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected148 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected149 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected150 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected151 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x13_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected144 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected145 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected146 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected147 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected148 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected149 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected150 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected151 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x14_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected152 | monroe_ionphoton_rtio_core_outputs_selected153) | monroe_ionphoton_rtio_core_outputs_selected154) | monroe_ionphoton_rtio_core_outputs_selected155) | monroe_ionphoton_rtio_core_outputs_selected156) | monroe_ionphoton_rtio_core_outputs_selected157) | monroe_ionphoton_rtio_core_outputs_selected158) | monroe_ionphoton_rtio_core_outputs_selected159);
	output_8x14_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected152 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected153 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected154 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected155 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected156 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected157 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected158 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected159 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x14_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected152 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected153 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected154 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected155 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected156 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected157 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected158 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected159 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x15_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected160 | monroe_ionphoton_rtio_core_outputs_selected161) | monroe_ionphoton_rtio_core_outputs_selected162) | monroe_ionphoton_rtio_core_outputs_selected163) | monroe_ionphoton_rtio_core_outputs_selected164) | monroe_ionphoton_rtio_core_outputs_selected165) | monroe_ionphoton_rtio_core_outputs_selected166) | monroe_ionphoton_rtio_core_outputs_selected167);
	output_8x15_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected160 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected161 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected162 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected163 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected164 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected165 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected166 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected167 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x15_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected160 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected161 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected162 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected163 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected164 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected165 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected166 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected167 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x16_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected168 | monroe_ionphoton_rtio_core_outputs_selected169) | monroe_ionphoton_rtio_core_outputs_selected170) | monroe_ionphoton_rtio_core_outputs_selected171) | monroe_ionphoton_rtio_core_outputs_selected172) | monroe_ionphoton_rtio_core_outputs_selected173) | monroe_ionphoton_rtio_core_outputs_selected174) | monroe_ionphoton_rtio_core_outputs_selected175);
	output_8x16_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected168 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected169 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected170 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected171 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected172 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected173 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected174 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected175 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x16_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected168 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected169 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected170 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected171 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected172 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected173 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected174 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected175 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	spimaster1_ointerface1_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected176 | monroe_ionphoton_rtio_core_outputs_selected177) | monroe_ionphoton_rtio_core_outputs_selected178) | monroe_ionphoton_rtio_core_outputs_selected179) | monroe_ionphoton_rtio_core_outputs_selected180) | monroe_ionphoton_rtio_core_outputs_selected181) | monroe_ionphoton_rtio_core_outputs_selected182) | monroe_ionphoton_rtio_core_outputs_selected183);
	spimaster1_ointerface1_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected176 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected177 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected178 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected179 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected180 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected181 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected182 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected183 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	spimaster1_ointerface1_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected176 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected177 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected178 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected179 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected180 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected181 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected182 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected183 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x17_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected184 | monroe_ionphoton_rtio_core_outputs_selected185) | monroe_ionphoton_rtio_core_outputs_selected186) | monroe_ionphoton_rtio_core_outputs_selected187) | monroe_ionphoton_rtio_core_outputs_selected188) | monroe_ionphoton_rtio_core_outputs_selected189) | monroe_ionphoton_rtio_core_outputs_selected190) | monroe_ionphoton_rtio_core_outputs_selected191);
	output_8x17_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected184 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected185 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected186 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected187 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected188 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected189 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected190 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected191 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x17_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected184 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected185 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected186 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected187 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected188 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected189 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected190 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected191 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x18_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected192 | monroe_ionphoton_rtio_core_outputs_selected193) | monroe_ionphoton_rtio_core_outputs_selected194) | monroe_ionphoton_rtio_core_outputs_selected195) | monroe_ionphoton_rtio_core_outputs_selected196) | monroe_ionphoton_rtio_core_outputs_selected197) | monroe_ionphoton_rtio_core_outputs_selected198) | monroe_ionphoton_rtio_core_outputs_selected199);
	output_8x18_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected192 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected193 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected194 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected195 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected196 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected197 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected198 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected199 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x18_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected192 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected193 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected194 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected195 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected196 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected197 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected198 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected199 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x19_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected200 | monroe_ionphoton_rtio_core_outputs_selected201) | monroe_ionphoton_rtio_core_outputs_selected202) | monroe_ionphoton_rtio_core_outputs_selected203) | monroe_ionphoton_rtio_core_outputs_selected204) | monroe_ionphoton_rtio_core_outputs_selected205) | monroe_ionphoton_rtio_core_outputs_selected206) | monroe_ionphoton_rtio_core_outputs_selected207);
	output_8x19_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected200 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected201 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected202 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected203 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected204 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected205 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected206 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected207 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x19_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected200 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected201 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected202 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected203 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected204 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected205 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected206 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected207 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x20_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected208 | monroe_ionphoton_rtio_core_outputs_selected209) | monroe_ionphoton_rtio_core_outputs_selected210) | monroe_ionphoton_rtio_core_outputs_selected211) | monroe_ionphoton_rtio_core_outputs_selected212) | monroe_ionphoton_rtio_core_outputs_selected213) | monroe_ionphoton_rtio_core_outputs_selected214) | monroe_ionphoton_rtio_core_outputs_selected215);
	output_8x20_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected208 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected209 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected210 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected211 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected212 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected213 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected214 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected215 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x20_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected208 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected209 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected210 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected211 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected212 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected213 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected214 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected215 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x21_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected216 | monroe_ionphoton_rtio_core_outputs_selected217) | monroe_ionphoton_rtio_core_outputs_selected218) | monroe_ionphoton_rtio_core_outputs_selected219) | monroe_ionphoton_rtio_core_outputs_selected220) | monroe_ionphoton_rtio_core_outputs_selected221) | monroe_ionphoton_rtio_core_outputs_selected222) | monroe_ionphoton_rtio_core_outputs_selected223);
	output_8x21_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected216 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected217 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected218 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected219 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected220 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected221 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected222 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected223 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x21_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected216 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected217 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected218 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected219 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected220 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected221 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected222 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected223 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	spimaster2_ointerface2_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected224 | monroe_ionphoton_rtio_core_outputs_selected225) | monroe_ionphoton_rtio_core_outputs_selected226) | monroe_ionphoton_rtio_core_outputs_selected227) | monroe_ionphoton_rtio_core_outputs_selected228) | monroe_ionphoton_rtio_core_outputs_selected229) | monroe_ionphoton_rtio_core_outputs_selected230) | monroe_ionphoton_rtio_core_outputs_selected231);
	spimaster2_ointerface2_address <= ((((((((monroe_ionphoton_rtio_core_outputs_selected224 ? monroe_ionphoton_rtio_core_outputs_record0_payload_address3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected225 ? monroe_ionphoton_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected226 ? monroe_ionphoton_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected227 ? monroe_ionphoton_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected228 ? monroe_ionphoton_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected229 ? monroe_ionphoton_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected230 ? monroe_ionphoton_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected231 ? monroe_ionphoton_rtio_core_outputs_record7_payload_address3 : 1'd0));
	spimaster2_ointerface2_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected224 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected225 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected226 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected227 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected228 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected229 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected230 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected231 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x22_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected232 | monroe_ionphoton_rtio_core_outputs_selected233) | monroe_ionphoton_rtio_core_outputs_selected234) | monroe_ionphoton_rtio_core_outputs_selected235) | monroe_ionphoton_rtio_core_outputs_selected236) | monroe_ionphoton_rtio_core_outputs_selected237) | monroe_ionphoton_rtio_core_outputs_selected238) | monroe_ionphoton_rtio_core_outputs_selected239);
	output_8x22_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected232 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected233 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected234 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected235 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected236 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected237 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected238 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected239 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x22_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected232 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected233 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected234 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected235 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected236 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected237 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected238 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected239 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x23_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected240 | monroe_ionphoton_rtio_core_outputs_selected241) | monroe_ionphoton_rtio_core_outputs_selected242) | monroe_ionphoton_rtio_core_outputs_selected243) | monroe_ionphoton_rtio_core_outputs_selected244) | monroe_ionphoton_rtio_core_outputs_selected245) | monroe_ionphoton_rtio_core_outputs_selected246) | monroe_ionphoton_rtio_core_outputs_selected247);
	output_8x23_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected240 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected241 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected242 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected243 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected244 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected245 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected246 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected247 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x23_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected240 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected241 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected242 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected243 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected244 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected245 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected246 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected247 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x24_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected248 | monroe_ionphoton_rtio_core_outputs_selected249) | monroe_ionphoton_rtio_core_outputs_selected250) | monroe_ionphoton_rtio_core_outputs_selected251) | monroe_ionphoton_rtio_core_outputs_selected252) | monroe_ionphoton_rtio_core_outputs_selected253) | monroe_ionphoton_rtio_core_outputs_selected254) | monroe_ionphoton_rtio_core_outputs_selected255);
	output_8x24_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected248 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected249 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected250 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected251 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected252 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected253 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected254 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected255 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x24_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected248 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected249 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected250 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected251 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected252 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected253 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected254 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected255 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x25_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected256 | monroe_ionphoton_rtio_core_outputs_selected257) | monroe_ionphoton_rtio_core_outputs_selected258) | monroe_ionphoton_rtio_core_outputs_selected259) | monroe_ionphoton_rtio_core_outputs_selected260) | monroe_ionphoton_rtio_core_outputs_selected261) | monroe_ionphoton_rtio_core_outputs_selected262) | monroe_ionphoton_rtio_core_outputs_selected263);
	output_8x25_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected256 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected257 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected258 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected259 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected260 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected261 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected262 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected263 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x25_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected256 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected257 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected258 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected259 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected260 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected261 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected262 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected263 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output_8x26_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected264 | monroe_ionphoton_rtio_core_outputs_selected265) | monroe_ionphoton_rtio_core_outputs_selected266) | monroe_ionphoton_rtio_core_outputs_selected267) | monroe_ionphoton_rtio_core_outputs_selected268) | monroe_ionphoton_rtio_core_outputs_selected269) | monroe_ionphoton_rtio_core_outputs_selected270) | monroe_ionphoton_rtio_core_outputs_selected271);
	output_8x26_fine_ts <= ((((((((monroe_ionphoton_rtio_core_outputs_selected264 ? monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected265 ? monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected266 ? monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected267 ? monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected268 ? monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected269 ? monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected270 ? monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected271 ? monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	output_8x26_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected264 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected265 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected266 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected267 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected268 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected269 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected270 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected271 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output0_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected272 | monroe_ionphoton_rtio_core_outputs_selected273) | monroe_ionphoton_rtio_core_outputs_selected274) | monroe_ionphoton_rtio_core_outputs_selected275) | monroe_ionphoton_rtio_core_outputs_selected276) | monroe_ionphoton_rtio_core_outputs_selected277) | monroe_ionphoton_rtio_core_outputs_selected278) | monroe_ionphoton_rtio_core_outputs_selected279);
	output0_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected272 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected273 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected274 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected275 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected276 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected277 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected278 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected279 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	output1_stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected280 | monroe_ionphoton_rtio_core_outputs_selected281) | monroe_ionphoton_rtio_core_outputs_selected282) | monroe_ionphoton_rtio_core_outputs_selected283) | monroe_ionphoton_rtio_core_outputs_selected284) | monroe_ionphoton_rtio_core_outputs_selected285) | monroe_ionphoton_rtio_core_outputs_selected286) | monroe_ionphoton_rtio_core_outputs_selected287);
	output1_data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected280 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected281 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected282 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected283 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected284 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected285 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected286 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected287 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	stb <= (((((((monroe_ionphoton_rtio_core_outputs_selected288 | monroe_ionphoton_rtio_core_outputs_selected289) | monroe_ionphoton_rtio_core_outputs_selected290) | monroe_ionphoton_rtio_core_outputs_selected291) | monroe_ionphoton_rtio_core_outputs_selected292) | monroe_ionphoton_rtio_core_outputs_selected293) | monroe_ionphoton_rtio_core_outputs_selected294) | monroe_ionphoton_rtio_core_outputs_selected295);
	data <= ((((((((monroe_ionphoton_rtio_core_outputs_selected288 ? monroe_ionphoton_rtio_core_outputs_record0_payload_data3 : 1'd0) | (monroe_ionphoton_rtio_core_outputs_selected289 ? monroe_ionphoton_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected290 ? monroe_ionphoton_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected291 ? monroe_ionphoton_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected292 ? monroe_ionphoton_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected293 ? monroe_ionphoton_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected294 ? monroe_ionphoton_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (monroe_ionphoton_rtio_core_outputs_selected295 ? monroe_ionphoton_rtio_core_outputs_record7_payload_data3 : 1'd0));
	monroe_ionphoton_rtio_core_outputs_busy <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_busy_channel <= 1'd0;
	monroe_ionphoton_rtio_core_outputs_stb_r0 <= (monroe_ionphoton_rtio_core_outputs_record0_valid1 & (~monroe_ionphoton_rtio_core_outputs_record0_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r0 <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r0 & sync_basiclowerer_array_muxed0)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r0;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r1 <= (monroe_ionphoton_rtio_core_outputs_record1_valid1 & (~monroe_ionphoton_rtio_core_outputs_record1_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r1 <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r1 & sync_basiclowerer_array_muxed1)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r1;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r2 <= (monroe_ionphoton_rtio_core_outputs_record2_valid1 & (~monroe_ionphoton_rtio_core_outputs_record2_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r2 <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r2 & sync_basiclowerer_array_muxed2)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r2;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r3 <= (monroe_ionphoton_rtio_core_outputs_record3_valid1 & (~monroe_ionphoton_rtio_core_outputs_record3_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r3 <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r3 & sync_basiclowerer_array_muxed3)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r3;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r4 <= (monroe_ionphoton_rtio_core_outputs_record4_valid1 & (~monroe_ionphoton_rtio_core_outputs_record4_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r4 <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r4 & sync_basiclowerer_array_muxed4)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r4;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r5 <= (monroe_ionphoton_rtio_core_outputs_record5_valid1 & (~monroe_ionphoton_rtio_core_outputs_record5_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r5 <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r5 & sync_basiclowerer_array_muxed5)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r5;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r6 <= (monroe_ionphoton_rtio_core_outputs_record6_valid1 & (~monroe_ionphoton_rtio_core_outputs_record6_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r6 <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r6 & sync_basiclowerer_array_muxed6)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r6;
	end
	monroe_ionphoton_rtio_core_outputs_stb_r7 <= (monroe_ionphoton_rtio_core_outputs_record7_valid1 & (~monroe_ionphoton_rtio_core_outputs_record7_collision));
	monroe_ionphoton_rtio_core_outputs_channel_r7 <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel3;
	if ((monroe_ionphoton_rtio_core_outputs_stb_r7 & sync_basiclowerer_array_muxed7)) begin
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_busy_channel <= monroe_ionphoton_rtio_core_outputs_channel_r7;
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record0_valid0), monroe_ionphoton_rtio_core_outputs_record0_payload_channel2} == {(~monroe_ionphoton_rtio_core_outputs_record1_valid0), monroe_ionphoton_rtio_core_outputs_record1_payload_channel2})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record0_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record0_seqn2[11]) & (monroe_ionphoton_rtio_core_outputs_record1_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record1_seqn2[11])) & (monroe_ionphoton_rtio_core_outputs_record0_seqn2[11] != monroe_ionphoton_rtio_core_outputs_record1_seqn2[11])) ? monroe_ionphoton_rtio_core_outputs_record0_seqn2[11] : (monroe_ionphoton_rtio_core_outputs_record0_seqn2 < monroe_ionphoton_rtio_core_outputs_record1_seqn2))) begin
			monroe_ionphoton_rtio_core_outputs_record0_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_valid0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_seqn2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_valid0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_seqn2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record0_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_valid0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_seqn2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_valid0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_seqn2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_payload_data2;
		end
		monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference0;
		monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record0_valid0), monroe_ionphoton_rtio_core_outputs_record0_payload_channel2} < {(~monroe_ionphoton_rtio_core_outputs_record1_valid0), monroe_ionphoton_rtio_core_outputs_record1_payload_channel2})) begin
			monroe_ionphoton_rtio_core_outputs_record0_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_valid0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_seqn2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_valid0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_seqn2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record0_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_valid0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_seqn2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_valid0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_seqn2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_payload_data2;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record2_valid0), monroe_ionphoton_rtio_core_outputs_record2_payload_channel2} == {(~monroe_ionphoton_rtio_core_outputs_record3_valid0), monroe_ionphoton_rtio_core_outputs_record3_payload_channel2})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record2_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record2_seqn2[11]) & (monroe_ionphoton_rtio_core_outputs_record3_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record3_seqn2[11])) & (monroe_ionphoton_rtio_core_outputs_record2_seqn2[11] != monroe_ionphoton_rtio_core_outputs_record3_seqn2[11])) ? monroe_ionphoton_rtio_core_outputs_record2_seqn2[11] : (monroe_ionphoton_rtio_core_outputs_record2_seqn2 < monroe_ionphoton_rtio_core_outputs_record3_seqn2))) begin
			monroe_ionphoton_rtio_core_outputs_record2_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_valid0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_seqn2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_valid0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_seqn2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record2_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_valid0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_seqn2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_valid0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_seqn2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_payload_data2;
		end
		monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference1;
		monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record2_valid0), monroe_ionphoton_rtio_core_outputs_record2_payload_channel2} < {(~monroe_ionphoton_rtio_core_outputs_record3_valid0), monroe_ionphoton_rtio_core_outputs_record3_payload_channel2})) begin
			monroe_ionphoton_rtio_core_outputs_record2_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_valid0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_seqn2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_valid0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_seqn2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record2_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_valid0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_seqn2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_valid0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_seqn2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_payload_data2;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record4_valid0), monroe_ionphoton_rtio_core_outputs_record4_payload_channel2} == {(~monroe_ionphoton_rtio_core_outputs_record5_valid0), monroe_ionphoton_rtio_core_outputs_record5_payload_channel2})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record4_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record4_seqn2[11]) & (monroe_ionphoton_rtio_core_outputs_record5_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record5_seqn2[11])) & (monroe_ionphoton_rtio_core_outputs_record4_seqn2[11] != monroe_ionphoton_rtio_core_outputs_record5_seqn2[11])) ? monroe_ionphoton_rtio_core_outputs_record4_seqn2[11] : (monroe_ionphoton_rtio_core_outputs_record4_seqn2 < monroe_ionphoton_rtio_core_outputs_record5_seqn2))) begin
			monroe_ionphoton_rtio_core_outputs_record4_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_valid0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_seqn2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_valid0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_seqn2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record4_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_valid0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_seqn2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_valid0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_seqn2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_payload_data2;
		end
		monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference2;
		monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record4_valid0), monroe_ionphoton_rtio_core_outputs_record4_payload_channel2} < {(~monroe_ionphoton_rtio_core_outputs_record5_valid0), monroe_ionphoton_rtio_core_outputs_record5_payload_channel2})) begin
			monroe_ionphoton_rtio_core_outputs_record4_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_valid0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_seqn2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_valid0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_seqn2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record4_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_valid0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_seqn2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_valid0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_seqn2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_payload_data2;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record6_valid0), monroe_ionphoton_rtio_core_outputs_record6_payload_channel2} == {(~monroe_ionphoton_rtio_core_outputs_record7_valid0), monroe_ionphoton_rtio_core_outputs_record7_payload_channel2})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record6_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record6_seqn2[11]) & (monroe_ionphoton_rtio_core_outputs_record7_seqn2[10] == monroe_ionphoton_rtio_core_outputs_record7_seqn2[11])) & (monroe_ionphoton_rtio_core_outputs_record6_seqn2[11] != monroe_ionphoton_rtio_core_outputs_record7_seqn2[11])) ? monroe_ionphoton_rtio_core_outputs_record6_seqn2[11] : (monroe_ionphoton_rtio_core_outputs_record6_seqn2 < monroe_ionphoton_rtio_core_outputs_record7_seqn2))) begin
			monroe_ionphoton_rtio_core_outputs_record6_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_valid0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_seqn2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_valid0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_seqn2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record6_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_valid0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_seqn2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_valid0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_seqn2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_payload_data2;
		end
		monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference3;
		monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record6_valid0), monroe_ionphoton_rtio_core_outputs_record6_payload_channel2} < {(~monroe_ionphoton_rtio_core_outputs_record7_valid0), monroe_ionphoton_rtio_core_outputs_record7_payload_channel2})) begin
			monroe_ionphoton_rtio_core_outputs_record6_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_valid0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_seqn2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_valid0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_seqn2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_payload_data2;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record6_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_valid0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_seqn2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_payload_data2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_valid0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_seqn2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_payload_channel2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_payload_fine_ts0;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_payload_address2;
			monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_payload_data2;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record0_rec_valid), monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record2_rec_valid), monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record0_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record0_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record2_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record2_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record0_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record2_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record0_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record0_rec_seqn < monroe_ionphoton_rtio_core_outputs_record2_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record8_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record8_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record10_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record8_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record8_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record10_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference4;
		monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record0_rec_valid), monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record2_rec_valid), monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record8_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record8_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record10_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record8_rec_valid <= monroe_ionphoton_rtio_core_outputs_record2_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record8_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record2_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record2_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record2_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= monroe_ionphoton_rtio_core_outputs_record0_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record10_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record0_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record0_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record0_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record1_rec_valid), monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record3_rec_valid), monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record1_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record1_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record3_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record3_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record1_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record3_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record1_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record1_rec_seqn < monroe_ionphoton_rtio_core_outputs_record3_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record9_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record9_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record11_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record9_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record9_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record11_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference5;
		monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record1_rec_valid), monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record3_rec_valid), monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record9_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record9_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record11_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record9_rec_valid <= monroe_ionphoton_rtio_core_outputs_record3_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record9_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record3_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record3_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record3_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= monroe_ionphoton_rtio_core_outputs_record1_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record11_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record1_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record1_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record1_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record4_rec_valid), monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record6_rec_valid), monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record4_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record4_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record6_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record6_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record4_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record6_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record4_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record4_rec_seqn < monroe_ionphoton_rtio_core_outputs_record6_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record12_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record12_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record14_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record12_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record12_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record14_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference6;
		monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record4_rec_valid), monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record6_rec_valid), monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record12_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record12_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record14_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record12_rec_valid <= monroe_ionphoton_rtio_core_outputs_record6_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record12_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record6_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record6_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record6_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= monroe_ionphoton_rtio_core_outputs_record4_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record14_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record4_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record4_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record4_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record5_rec_valid), monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record7_rec_valid), monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record5_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record5_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record7_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record7_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record5_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record7_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record5_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record5_rec_seqn < monroe_ionphoton_rtio_core_outputs_record7_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record13_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record13_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record15_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record13_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record13_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record15_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference7;
		monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record5_rec_valid), monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record7_rec_valid), monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record13_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record13_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record15_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record13_rec_valid <= monroe_ionphoton_rtio_core_outputs_record7_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record13_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record7_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record7_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record7_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= monroe_ionphoton_rtio_core_outputs_record5_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record15_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record5_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record5_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record5_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record9_rec_valid), monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record10_rec_valid), monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record9_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record9_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record10_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record10_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record9_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record10_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record9_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record9_rec_seqn < monroe_ionphoton_rtio_core_outputs_record10_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record17_rec_valid <= monroe_ionphoton_rtio_core_outputs_record10_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record17_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record10_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= monroe_ionphoton_rtio_core_outputs_record9_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record18_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record9_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record17_rec_valid <= monroe_ionphoton_rtio_core_outputs_record9_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record17_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record9_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= monroe_ionphoton_rtio_core_outputs_record10_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record18_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record10_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference8;
		monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record9_rec_valid), monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record10_rec_valid), monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record17_rec_valid <= monroe_ionphoton_rtio_core_outputs_record9_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record17_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record9_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= monroe_ionphoton_rtio_core_outputs_record10_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record18_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record10_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record17_rec_valid <= monroe_ionphoton_rtio_core_outputs_record10_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record17_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record10_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record10_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record10_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= monroe_ionphoton_rtio_core_outputs_record9_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record18_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record9_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record9_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record9_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record13_rec_valid), monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record14_rec_valid), monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record13_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record13_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record14_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record14_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record13_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record14_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record13_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record13_rec_seqn < monroe_ionphoton_rtio_core_outputs_record14_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record21_rec_valid <= monroe_ionphoton_rtio_core_outputs_record14_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record21_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record14_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= monroe_ionphoton_rtio_core_outputs_record13_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record22_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record13_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record21_rec_valid <= monroe_ionphoton_rtio_core_outputs_record13_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record21_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record13_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= monroe_ionphoton_rtio_core_outputs_record14_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record22_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record14_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference9;
		monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record13_rec_valid), monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record14_rec_valid), monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record21_rec_valid <= monroe_ionphoton_rtio_core_outputs_record13_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record21_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record13_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= monroe_ionphoton_rtio_core_outputs_record14_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record22_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record14_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record21_rec_valid <= monroe_ionphoton_rtio_core_outputs_record14_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record21_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record14_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record14_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record14_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= monroe_ionphoton_rtio_core_outputs_record13_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record22_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record13_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record13_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record13_rec_payload_data;
		end
	end
	monroe_ionphoton_rtio_core_outputs_record16_rec_valid <= monroe_ionphoton_rtio_core_outputs_record8_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record16_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record8_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record8_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record8_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record8_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record8_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record8_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record8_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record19_rec_valid <= monroe_ionphoton_rtio_core_outputs_record11_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record19_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record11_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record11_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record11_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record11_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record11_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record11_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record11_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record20_rec_valid <= monroe_ionphoton_rtio_core_outputs_record12_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record20_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record12_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record12_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record12_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record12_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record12_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record12_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record12_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record23_rec_valid <= monroe_ionphoton_rtio_core_outputs_record15_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record23_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record15_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record15_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record15_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record15_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record15_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record15_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record15_rec_payload_data;
	if (({(~monroe_ionphoton_rtio_core_outputs_record16_rec_valid), monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record20_rec_valid), monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record16_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record16_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record20_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record20_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record16_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record20_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record16_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record16_rec_seqn < monroe_ionphoton_rtio_core_outputs_record20_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record24_rec_valid <= monroe_ionphoton_rtio_core_outputs_record20_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record24_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record20_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= monroe_ionphoton_rtio_core_outputs_record16_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record28_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record16_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record24_rec_valid <= monroe_ionphoton_rtio_core_outputs_record16_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record24_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record16_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= monroe_ionphoton_rtio_core_outputs_record20_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record28_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record20_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference10;
		monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record16_rec_valid), monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record20_rec_valid), monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record24_rec_valid <= monroe_ionphoton_rtio_core_outputs_record16_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record24_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record16_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= monroe_ionphoton_rtio_core_outputs_record20_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record28_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record20_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record24_rec_valid <= monroe_ionphoton_rtio_core_outputs_record20_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record24_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record20_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record20_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record20_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= monroe_ionphoton_rtio_core_outputs_record16_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record28_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record16_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record16_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record16_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record17_rec_valid), monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record21_rec_valid), monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record17_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record17_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record21_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record21_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record17_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record21_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record17_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record17_rec_seqn < monroe_ionphoton_rtio_core_outputs_record21_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record25_rec_valid <= monroe_ionphoton_rtio_core_outputs_record21_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record25_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record21_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= monroe_ionphoton_rtio_core_outputs_record17_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record29_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record17_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record25_rec_valid <= monroe_ionphoton_rtio_core_outputs_record17_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record25_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record17_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= monroe_ionphoton_rtio_core_outputs_record21_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record29_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record21_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference11;
		monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record17_rec_valid), monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record21_rec_valid), monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record25_rec_valid <= monroe_ionphoton_rtio_core_outputs_record17_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record25_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record17_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= monroe_ionphoton_rtio_core_outputs_record21_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record29_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record21_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record25_rec_valid <= monroe_ionphoton_rtio_core_outputs_record21_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record25_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record21_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record21_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record21_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= monroe_ionphoton_rtio_core_outputs_record17_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record29_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record17_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record17_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record17_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record18_rec_valid), monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record22_rec_valid), monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record18_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record18_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record22_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record22_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record18_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record22_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record18_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record18_rec_seqn < monroe_ionphoton_rtio_core_outputs_record22_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record26_rec_valid <= monroe_ionphoton_rtio_core_outputs_record22_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record26_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record22_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= monroe_ionphoton_rtio_core_outputs_record18_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record30_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record18_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record26_rec_valid <= monroe_ionphoton_rtio_core_outputs_record18_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record26_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record18_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= monroe_ionphoton_rtio_core_outputs_record22_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record30_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record22_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference12;
		monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record18_rec_valid), monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record22_rec_valid), monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record26_rec_valid <= monroe_ionphoton_rtio_core_outputs_record18_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record26_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record18_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= monroe_ionphoton_rtio_core_outputs_record22_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record30_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record22_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record26_rec_valid <= monroe_ionphoton_rtio_core_outputs_record22_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record26_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record22_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record22_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record22_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= monroe_ionphoton_rtio_core_outputs_record18_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record30_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record18_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record18_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record18_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record19_rec_valid), monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record23_rec_valid), monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record19_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record19_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record23_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record23_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record19_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record23_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record19_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record19_rec_seqn < monroe_ionphoton_rtio_core_outputs_record23_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record27_rec_valid <= monroe_ionphoton_rtio_core_outputs_record23_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record27_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record23_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= monroe_ionphoton_rtio_core_outputs_record19_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record31_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record19_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record27_rec_valid <= monroe_ionphoton_rtio_core_outputs_record19_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record27_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record19_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= monroe_ionphoton_rtio_core_outputs_record23_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record31_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record23_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference13;
		monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record19_rec_valid), monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record23_rec_valid), monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record27_rec_valid <= monroe_ionphoton_rtio_core_outputs_record19_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record27_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record19_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= monroe_ionphoton_rtio_core_outputs_record23_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record31_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record23_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record27_rec_valid <= monroe_ionphoton_rtio_core_outputs_record23_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record27_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record23_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record23_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record23_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= monroe_ionphoton_rtio_core_outputs_record19_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record31_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record19_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record19_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record19_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record26_rec_valid), monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record28_rec_valid), monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record26_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record26_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record28_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record28_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record26_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record28_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record26_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record26_rec_seqn < monroe_ionphoton_rtio_core_outputs_record28_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record34_rec_valid <= monroe_ionphoton_rtio_core_outputs_record28_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record34_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record28_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= monroe_ionphoton_rtio_core_outputs_record26_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record36_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record26_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record34_rec_valid <= monroe_ionphoton_rtio_core_outputs_record26_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record34_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record26_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= monroe_ionphoton_rtio_core_outputs_record28_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record36_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record28_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference14;
		monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record26_rec_valid), monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record28_rec_valid), monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record34_rec_valid <= monroe_ionphoton_rtio_core_outputs_record26_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record34_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record26_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= monroe_ionphoton_rtio_core_outputs_record28_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record36_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record28_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record34_rec_valid <= monroe_ionphoton_rtio_core_outputs_record28_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record34_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record28_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record28_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record28_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= monroe_ionphoton_rtio_core_outputs_record26_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record36_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record26_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record26_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record26_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record27_rec_valid), monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record29_rec_valid), monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record27_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record27_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record29_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record29_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record27_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record29_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record27_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record27_rec_seqn < monroe_ionphoton_rtio_core_outputs_record29_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record35_rec_valid <= monroe_ionphoton_rtio_core_outputs_record29_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record35_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record29_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= monroe_ionphoton_rtio_core_outputs_record27_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record37_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record27_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record35_rec_valid <= monroe_ionphoton_rtio_core_outputs_record27_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record35_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record27_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= monroe_ionphoton_rtio_core_outputs_record29_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record37_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record29_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference15;
		monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record27_rec_valid), monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record29_rec_valid), monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record35_rec_valid <= monroe_ionphoton_rtio_core_outputs_record27_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record35_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record27_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= monroe_ionphoton_rtio_core_outputs_record29_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record37_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record29_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record35_rec_valid <= monroe_ionphoton_rtio_core_outputs_record29_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record35_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record29_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record29_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record29_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= monroe_ionphoton_rtio_core_outputs_record27_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record37_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record27_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record27_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record27_rec_payload_data;
		end
	end
	monroe_ionphoton_rtio_core_outputs_record32_rec_valid <= monroe_ionphoton_rtio_core_outputs_record24_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record32_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record24_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record32_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record24_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record32_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record24_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record32_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record24_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record32_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record24_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record32_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record24_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record32_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record24_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record33_rec_valid <= monroe_ionphoton_rtio_core_outputs_record25_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record33_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record25_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record25_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record25_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record25_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record25_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record25_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record25_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record38_rec_valid <= monroe_ionphoton_rtio_core_outputs_record30_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record38_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record30_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record30_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record30_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record30_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record30_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record30_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record30_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record39_rec_valid <= monroe_ionphoton_rtio_core_outputs_record31_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record39_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record31_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record39_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record31_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record39_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record31_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record39_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record31_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record39_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record31_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record39_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record31_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record39_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record31_rec_payload_data;
	if (({(~monroe_ionphoton_rtio_core_outputs_record33_rec_valid), monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record34_rec_valid), monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record33_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record33_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record34_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record34_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record33_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record34_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record33_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record33_rec_seqn < monroe_ionphoton_rtio_core_outputs_record34_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record41_rec_valid <= monroe_ionphoton_rtio_core_outputs_record34_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record41_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record34_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= monroe_ionphoton_rtio_core_outputs_record33_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record42_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record33_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record41_rec_valid <= monroe_ionphoton_rtio_core_outputs_record33_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record41_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record33_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= monroe_ionphoton_rtio_core_outputs_record34_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record42_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record34_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference16;
		monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record33_rec_valid), monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record34_rec_valid), monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record41_rec_valid <= monroe_ionphoton_rtio_core_outputs_record33_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record41_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record33_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= monroe_ionphoton_rtio_core_outputs_record34_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record42_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record34_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record41_rec_valid <= monroe_ionphoton_rtio_core_outputs_record34_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record41_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record34_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record41_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record34_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record41_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record34_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= monroe_ionphoton_rtio_core_outputs_record33_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record42_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record33_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record42_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record33_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record42_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record33_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record35_rec_valid), monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record36_rec_valid), monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record35_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record35_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record36_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record36_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record35_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record36_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record35_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record35_rec_seqn < monroe_ionphoton_rtio_core_outputs_record36_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record43_rec_valid <= monroe_ionphoton_rtio_core_outputs_record36_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record43_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record36_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= monroe_ionphoton_rtio_core_outputs_record35_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record44_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record35_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record43_rec_valid <= monroe_ionphoton_rtio_core_outputs_record35_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record43_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record35_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= monroe_ionphoton_rtio_core_outputs_record36_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record44_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record36_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference17;
		monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record35_rec_valid), monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record36_rec_valid), monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record43_rec_valid <= monroe_ionphoton_rtio_core_outputs_record35_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record43_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record35_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= monroe_ionphoton_rtio_core_outputs_record36_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record44_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record36_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record43_rec_valid <= monroe_ionphoton_rtio_core_outputs_record36_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record43_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record36_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record43_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record36_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record43_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record36_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= monroe_ionphoton_rtio_core_outputs_record35_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record44_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record35_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record44_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record35_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record44_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record35_rec_payload_data;
		end
	end
	if (({(~monroe_ionphoton_rtio_core_outputs_record37_rec_valid), monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel} == {(~monroe_ionphoton_rtio_core_outputs_record38_rec_valid), monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel})) begin
		if (((((monroe_ionphoton_rtio_core_outputs_record37_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record37_rec_seqn[11]) & (monroe_ionphoton_rtio_core_outputs_record38_rec_seqn[10] == monroe_ionphoton_rtio_core_outputs_record38_rec_seqn[11])) & (monroe_ionphoton_rtio_core_outputs_record37_rec_seqn[11] != monroe_ionphoton_rtio_core_outputs_record38_rec_seqn[11])) ? monroe_ionphoton_rtio_core_outputs_record37_rec_seqn[11] : (monroe_ionphoton_rtio_core_outputs_record37_rec_seqn < monroe_ionphoton_rtio_core_outputs_record38_rec_seqn))) begin
			monroe_ionphoton_rtio_core_outputs_record45_rec_valid <= monroe_ionphoton_rtio_core_outputs_record38_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record45_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record38_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= monroe_ionphoton_rtio_core_outputs_record37_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record46_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record37_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record45_rec_valid <= monroe_ionphoton_rtio_core_outputs_record37_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record45_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record37_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= monroe_ionphoton_rtio_core_outputs_record38_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record46_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record38_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data;
		end
		monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_nondata_difference18;
		monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= 1'd0;
	end else begin
		if (({(~monroe_ionphoton_rtio_core_outputs_record37_rec_valid), monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel} < {(~monroe_ionphoton_rtio_core_outputs_record38_rec_valid), monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel})) begin
			monroe_ionphoton_rtio_core_outputs_record45_rec_valid <= monroe_ionphoton_rtio_core_outputs_record37_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record45_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record37_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= monroe_ionphoton_rtio_core_outputs_record38_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record46_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record38_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data;
		end else begin
			monroe_ionphoton_rtio_core_outputs_record45_rec_valid <= monroe_ionphoton_rtio_core_outputs_record38_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record45_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record38_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record45_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record38_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record45_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record38_rec_payload_data;
			monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= monroe_ionphoton_rtio_core_outputs_record37_rec_valid;
			monroe_ionphoton_rtio_core_outputs_record46_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record37_rec_seqn;
			monroe_ionphoton_rtio_core_outputs_record46_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record37_rec_nondata_replace_occured;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_channel;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_fine_ts;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_address;
			monroe_ionphoton_rtio_core_outputs_record46_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record37_rec_payload_data;
		end
	end
	monroe_ionphoton_rtio_core_outputs_record40_rec_valid <= monroe_ionphoton_rtio_core_outputs_record32_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record40_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record32_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record40_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record32_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record40_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record32_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record40_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record32_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record40_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record32_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record40_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record32_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record40_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record32_rec_payload_data;
	monroe_ionphoton_rtio_core_outputs_record47_rec_valid <= monroe_ionphoton_rtio_core_outputs_record39_rec_valid;
	monroe_ionphoton_rtio_core_outputs_record47_rec_seqn <= monroe_ionphoton_rtio_core_outputs_record39_rec_seqn;
	monroe_ionphoton_rtio_core_outputs_record47_rec_replace_occured <= monroe_ionphoton_rtio_core_outputs_record39_rec_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record47_rec_nondata_replace_occured <= monroe_ionphoton_rtio_core_outputs_record39_rec_nondata_replace_occured;
	monroe_ionphoton_rtio_core_outputs_record47_rec_payload_channel <= monroe_ionphoton_rtio_core_outputs_record39_rec_payload_channel;
	monroe_ionphoton_rtio_core_outputs_record47_rec_payload_fine_ts <= monroe_ionphoton_rtio_core_outputs_record39_rec_payload_fine_ts;
	monroe_ionphoton_rtio_core_outputs_record47_rec_payload_address <= monroe_ionphoton_rtio_core_outputs_record39_rec_payload_address;
	monroe_ionphoton_rtio_core_outputs_record47_rec_payload_data <= monroe_ionphoton_rtio_core_outputs_record39_rec_payload_data;
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer0_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer0_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer1_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer1_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer2_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer2_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer3_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer3_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer4_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer4_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer5_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer5_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer6_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer6_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_o) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
	if (monroe_ionphoton_rtio_core_o_collision_sync_i) begin
		monroe_ionphoton_rtio_core_o_collision_sync_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_o) begin
		monroe_ionphoton_rtio_core_o_collision_sync_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_o_collision_sync_ps_i) begin
		monroe_ionphoton_rtio_core_o_collision_sync_bxfer_data <= monroe_ionphoton_rtio_core_o_collision_sync_data_i;
	end
	if (monroe_ionphoton_rtio_core_o_collision_sync_ps_i) begin
		monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_i <= (~monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_o;
	if (monroe_ionphoton_rtio_core_o_busy_sync_i) begin
		monroe_ionphoton_rtio_core_o_busy_sync_blind <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_o) begin
		monroe_ionphoton_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_o_busy_sync_ps_i) begin
		monroe_ionphoton_rtio_core_o_busy_sync_bxfer_data <= monroe_ionphoton_rtio_core_o_busy_sync_data_i;
	end
	if (monroe_ionphoton_rtio_core_o_busy_sync_ps_i) begin
		monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_i <= (~monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_i);
	end
	monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o_r <= monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_o;
	if (rio_rst) begin
		inout_8x0_inout_8x0_ointerface0_stb <= 1'd0;
		inout_8x0_inout_8x0_sensitivity <= 2'd0;
		inout_8x0_inout_8x0_sample <= 1'd0;
		inout_8x1_inout_8x1_ointerface1_stb <= 1'd0;
		inout_8x1_inout_8x1_sensitivity <= 2'd0;
		inout_8x1_inout_8x1_sample <= 1'd0;
		inout_8x2_inout_8x2_ointerface2_stb <= 1'd0;
		inout_8x2_inout_8x2_sensitivity <= 2'd0;
		inout_8x2_inout_8x2_sample <= 1'd0;
		inout_8x3_inout_8x3_ointerface3_stb <= 1'd0;
		inout_8x3_inout_8x3_sensitivity <= 2'd0;
		inout_8x3_inout_8x3_sample <= 1'd0;
		output_8x0_stb <= 1'd0;
		output_8x1_stb <= 1'd0;
		output_8x2_stb <= 1'd0;
		output_8x3_stb <= 1'd0;
		output_8x4_stb <= 1'd0;
		output_8x5_stb <= 1'd0;
		output_8x6_stb <= 1'd0;
		output_8x7_stb <= 1'd0;
		output_8x8_stb <= 1'd0;
		output_8x9_stb <= 1'd0;
		output_8x10_stb <= 1'd0;
		output_8x11_stb <= 1'd0;
		spimaster0_ointerface0_stb <= 1'd0;
		output_8x12_stb <= 1'd0;
		output_8x13_stb <= 1'd0;
		output_8x14_stb <= 1'd0;
		output_8x15_stb <= 1'd0;
		output_8x16_stb <= 1'd0;
		spimaster1_ointerface1_stb <= 1'd0;
		output_8x17_stb <= 1'd0;
		output_8x18_stb <= 1'd0;
		output_8x19_stb <= 1'd0;
		output_8x20_stb <= 1'd0;
		output_8x21_stb <= 1'd0;
		spimaster2_ointerface2_stb <= 1'd0;
		output_8x22_stb <= 1'd0;
		output_8x23_stb <= 1'd0;
		output_8x24_stb <= 1'd0;
		output_8x25_stb <= 1'd0;
		output_8x26_stb <= 1'd0;
		output0_stb <= 1'd0;
		output1_stb <= 1'd0;
		stb <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_readable <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record0_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record1_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record2_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record3_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record4_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record5_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record6_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_gates_record7_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_collision <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_busy <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record0_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record1_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record2_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record3_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record4_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record5_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record6_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record7_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record8_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record9_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record10_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record11_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record12_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record13_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record14_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record15_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record16_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record17_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record18_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record19_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record20_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record21_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record22_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record23_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record24_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record25_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record26_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record27_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record28_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record29_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record30_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record31_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record32_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record33_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record34_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record35_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record36_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record37_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record38_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record39_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record40_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record41_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record42_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record43_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record44_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record45_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record46_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record47_rec_valid <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record0_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record1_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record2_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record3_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record4_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record5_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record6_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_record7_valid1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r0 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r0 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r2 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r2 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r3 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r3 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r4 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r4 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r5 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r5 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r6 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r6 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_replace_occured_r7 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_nondata_replace_occured_r7 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r0 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r1 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r2 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r3 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r4 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r5 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r6 <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_stb_r7 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
		monroe_ionphoton_rtio_core_o_collision_sync_blind <= 1'd0;
		monroe_ionphoton_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	xilinxmultiregimpl17_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q;
	xilinxmultiregimpl17_regs1 <= xilinxmultiregimpl17_regs0;
	xilinxmultiregimpl19_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q;
	xilinxmultiregimpl19_regs1 <= xilinxmultiregimpl19_regs0;
	xilinxmultiregimpl21_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q;
	xilinxmultiregimpl21_regs1 <= xilinxmultiregimpl21_regs0;
	xilinxmultiregimpl23_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q;
	xilinxmultiregimpl23_regs1 <= xilinxmultiregimpl23_regs0;
	xilinxmultiregimpl25_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q;
	xilinxmultiregimpl25_regs1 <= xilinxmultiregimpl25_regs0;
	xilinxmultiregimpl27_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q;
	xilinxmultiregimpl27_regs1 <= xilinxmultiregimpl27_regs0;
	xilinxmultiregimpl29_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q;
	xilinxmultiregimpl29_regs1 <= xilinxmultiregimpl29_regs0;
	xilinxmultiregimpl31_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q;
	xilinxmultiregimpl31_regs1 <= xilinxmultiregimpl31_regs0;
	xilinxmultiregimpl34_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q;
	xilinxmultiregimpl34_regs1 <= xilinxmultiregimpl34_regs0;
	xilinxmultiregimpl36_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i;
	xilinxmultiregimpl36_regs1 <= xilinxmultiregimpl36_regs0;
	xilinxmultiregimpl38_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q;
	xilinxmultiregimpl38_regs1 <= xilinxmultiregimpl38_regs0;
	xilinxmultiregimpl40_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i;
	xilinxmultiregimpl40_regs1 <= xilinxmultiregimpl40_regs0;
	xilinxmultiregimpl42_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q;
	xilinxmultiregimpl42_regs1 <= xilinxmultiregimpl42_regs0;
	xilinxmultiregimpl44_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i;
	xilinxmultiregimpl44_regs1 <= xilinxmultiregimpl44_regs0;
	xilinxmultiregimpl46_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q;
	xilinxmultiregimpl46_regs1 <= xilinxmultiregimpl46_regs0;
	xilinxmultiregimpl48_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i;
	xilinxmultiregimpl48_regs1 <= xilinxmultiregimpl48_regs0;
	xilinxmultiregimpl50_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q;
	xilinxmultiregimpl50_regs1 <= xilinxmultiregimpl50_regs0;
	xilinxmultiregimpl52_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i;
	xilinxmultiregimpl52_regs1 <= xilinxmultiregimpl52_regs0;
	xilinxmultiregimpl54_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q;
	xilinxmultiregimpl54_regs1 <= xilinxmultiregimpl54_regs0;
	xilinxmultiregimpl56_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i;
	xilinxmultiregimpl56_regs1 <= xilinxmultiregimpl56_regs0;
	xilinxmultiregimpl58_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q;
	xilinxmultiregimpl58_regs1 <= xilinxmultiregimpl58_regs0;
	xilinxmultiregimpl60_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i;
	xilinxmultiregimpl60_regs1 <= xilinxmultiregimpl60_regs0;
	xilinxmultiregimpl62_regs0 <= monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_i;
	xilinxmultiregimpl62_regs1 <= xilinxmultiregimpl62_regs0;
	xilinxmultiregimpl65_regs0 <= monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_i;
	xilinxmultiregimpl65_regs1 <= xilinxmultiregimpl65_regs0;
	xilinxmultiregimpl104_regs0 <= monroe_ionphoton_inj_o_sys0;
	xilinxmultiregimpl104_regs1 <= xilinxmultiregimpl104_regs0;
	xilinxmultiregimpl105_regs0 <= monroe_ionphoton_inj_o_sys1;
	xilinxmultiregimpl105_regs1 <= xilinxmultiregimpl105_regs0;
	xilinxmultiregimpl106_regs0 <= monroe_ionphoton_inj_o_sys2;
	xilinxmultiregimpl106_regs1 <= xilinxmultiregimpl106_regs0;
	xilinxmultiregimpl107_regs0 <= monroe_ionphoton_inj_o_sys3;
	xilinxmultiregimpl107_regs1 <= xilinxmultiregimpl107_regs0;
	xilinxmultiregimpl108_regs0 <= monroe_ionphoton_inj_o_sys4;
	xilinxmultiregimpl108_regs1 <= xilinxmultiregimpl108_regs0;
	xilinxmultiregimpl109_regs0 <= monroe_ionphoton_inj_o_sys5;
	xilinxmultiregimpl109_regs1 <= xilinxmultiregimpl109_regs0;
	xilinxmultiregimpl110_regs0 <= monroe_ionphoton_inj_o_sys6;
	xilinxmultiregimpl110_regs1 <= xilinxmultiregimpl110_regs0;
	xilinxmultiregimpl111_regs0 <= monroe_ionphoton_inj_o_sys7;
	xilinxmultiregimpl111_regs1 <= xilinxmultiregimpl111_regs0;
	xilinxmultiregimpl112_regs0 <= monroe_ionphoton_inj_o_sys8;
	xilinxmultiregimpl112_regs1 <= xilinxmultiregimpl112_regs0;
	xilinxmultiregimpl113_regs0 <= monroe_ionphoton_inj_o_sys9;
	xilinxmultiregimpl113_regs1 <= xilinxmultiregimpl113_regs0;
	xilinxmultiregimpl114_regs0 <= monroe_ionphoton_inj_o_sys10;
	xilinxmultiregimpl114_regs1 <= xilinxmultiregimpl114_regs0;
	xilinxmultiregimpl115_regs0 <= monroe_ionphoton_inj_o_sys11;
	xilinxmultiregimpl115_regs1 <= xilinxmultiregimpl115_regs0;
	xilinxmultiregimpl116_regs0 <= monroe_ionphoton_inj_o_sys12;
	xilinxmultiregimpl116_regs1 <= xilinxmultiregimpl116_regs0;
	xilinxmultiregimpl117_regs0 <= monroe_ionphoton_inj_o_sys13;
	xilinxmultiregimpl117_regs1 <= xilinxmultiregimpl117_regs0;
	xilinxmultiregimpl118_regs0 <= monroe_ionphoton_inj_o_sys14;
	xilinxmultiregimpl118_regs1 <= xilinxmultiregimpl118_regs0;
	xilinxmultiregimpl119_regs0 <= monroe_ionphoton_inj_o_sys15;
	xilinxmultiregimpl119_regs1 <= xilinxmultiregimpl119_regs0;
	xilinxmultiregimpl120_regs0 <= monroe_ionphoton_inj_o_sys16;
	xilinxmultiregimpl120_regs1 <= xilinxmultiregimpl120_regs0;
	xilinxmultiregimpl121_regs0 <= monroe_ionphoton_inj_o_sys17;
	xilinxmultiregimpl121_regs1 <= xilinxmultiregimpl121_regs0;
	xilinxmultiregimpl122_regs0 <= monroe_ionphoton_inj_o_sys18;
	xilinxmultiregimpl122_regs1 <= xilinxmultiregimpl122_regs0;
	xilinxmultiregimpl123_regs0 <= monroe_ionphoton_inj_o_sys19;
	xilinxmultiregimpl123_regs1 <= xilinxmultiregimpl123_regs0;
	xilinxmultiregimpl124_regs0 <= monroe_ionphoton_inj_o_sys20;
	xilinxmultiregimpl124_regs1 <= xilinxmultiregimpl124_regs0;
	xilinxmultiregimpl125_regs0 <= monroe_ionphoton_inj_o_sys21;
	xilinxmultiregimpl125_regs1 <= xilinxmultiregimpl125_regs0;
	xilinxmultiregimpl126_regs0 <= monroe_ionphoton_inj_o_sys22;
	xilinxmultiregimpl126_regs1 <= xilinxmultiregimpl126_regs0;
	xilinxmultiregimpl127_regs0 <= monroe_ionphoton_inj_o_sys23;
	xilinxmultiregimpl127_regs1 <= xilinxmultiregimpl127_regs0;
	xilinxmultiregimpl128_regs0 <= monroe_ionphoton_inj_o_sys24;
	xilinxmultiregimpl128_regs1 <= xilinxmultiregimpl128_regs0;
	xilinxmultiregimpl129_regs0 <= monroe_ionphoton_inj_o_sys25;
	xilinxmultiregimpl129_regs1 <= xilinxmultiregimpl129_regs0;
	xilinxmultiregimpl130_regs0 <= monroe_ionphoton_inj_o_sys26;
	xilinxmultiregimpl130_regs1 <= xilinxmultiregimpl130_regs0;
	xilinxmultiregimpl131_regs0 <= monroe_ionphoton_inj_o_sys27;
	xilinxmultiregimpl131_regs1 <= xilinxmultiregimpl131_regs0;
	xilinxmultiregimpl132_regs0 <= monroe_ionphoton_inj_o_sys28;
	xilinxmultiregimpl132_regs1 <= xilinxmultiregimpl132_regs0;
	xilinxmultiregimpl133_regs0 <= monroe_ionphoton_inj_o_sys29;
	xilinxmultiregimpl133_regs1 <= xilinxmultiregimpl133_regs0;
	xilinxmultiregimpl134_regs0 <= monroe_ionphoton_inj_o_sys30;
	xilinxmultiregimpl134_regs1 <= xilinxmultiregimpl134_regs0;
	xilinxmultiregimpl135_regs0 <= monroe_ionphoton_inj_o_sys31;
	xilinxmultiregimpl135_regs1 <= xilinxmultiregimpl135_regs0;
	xilinxmultiregimpl136_regs0 <= monroe_ionphoton_inj_o_sys32;
	xilinxmultiregimpl136_regs1 <= xilinxmultiregimpl136_regs0;
	xilinxmultiregimpl137_regs0 <= monroe_ionphoton_inj_o_sys33;
	xilinxmultiregimpl137_regs1 <= xilinxmultiregimpl137_regs0;
	xilinxmultiregimpl138_regs0 <= monroe_ionphoton_inj_o_sys34;
	xilinxmultiregimpl138_regs1 <= xilinxmultiregimpl138_regs0;
	xilinxmultiregimpl139_regs0 <= monroe_ionphoton_inj_o_sys35;
	xilinxmultiregimpl139_regs1 <= xilinxmultiregimpl139_regs0;
	xilinxmultiregimpl140_regs0 <= monroe_ionphoton_inj_o_sys36;
	xilinxmultiregimpl140_regs1 <= xilinxmultiregimpl140_regs0;
	xilinxmultiregimpl141_regs0 <= monroe_ionphoton_inj_o_sys37;
	xilinxmultiregimpl141_regs1 <= xilinxmultiregimpl141_regs0;
	xilinxmultiregimpl142_regs0 <= monroe_ionphoton_inj_o_sys38;
	xilinxmultiregimpl142_regs1 <= xilinxmultiregimpl142_regs0;
	xilinxmultiregimpl143_regs0 <= monroe_ionphoton_inj_o_sys39;
	xilinxmultiregimpl143_regs1 <= xilinxmultiregimpl143_regs0;
	xilinxmultiregimpl144_regs0 <= monroe_ionphoton_inj_o_sys40;
	xilinxmultiregimpl144_regs1 <= xilinxmultiregimpl144_regs0;
	xilinxmultiregimpl145_regs0 <= monroe_ionphoton_inj_o_sys41;
	xilinxmultiregimpl145_regs1 <= xilinxmultiregimpl145_regs0;
	xilinxmultiregimpl146_regs0 <= monroe_ionphoton_inj_o_sys42;
	xilinxmultiregimpl146_regs1 <= xilinxmultiregimpl146_regs0;
	xilinxmultiregimpl147_regs0 <= monroe_ionphoton_inj_o_sys43;
	xilinxmultiregimpl147_regs1 <= xilinxmultiregimpl147_regs0;
	xilinxmultiregimpl148_regs0 <= monroe_ionphoton_inj_o_sys44;
	xilinxmultiregimpl148_regs1 <= xilinxmultiregimpl148_regs0;
	xilinxmultiregimpl149_regs0 <= monroe_ionphoton_inj_o_sys45;
	xilinxmultiregimpl149_regs1 <= xilinxmultiregimpl149_regs0;
	xilinxmultiregimpl150_regs0 <= monroe_ionphoton_inj_o_sys46;
	xilinxmultiregimpl150_regs1 <= xilinxmultiregimpl150_regs0;
	xilinxmultiregimpl151_regs0 <= monroe_ionphoton_inj_o_sys47;
	xilinxmultiregimpl151_regs1 <= xilinxmultiregimpl151_regs0;
	xilinxmultiregimpl152_regs0 <= monroe_ionphoton_inj_o_sys48;
	xilinxmultiregimpl152_regs1 <= xilinxmultiregimpl152_regs0;
	xilinxmultiregimpl153_regs0 <= monroe_ionphoton_inj_o_sys49;
	xilinxmultiregimpl153_regs1 <= xilinxmultiregimpl153_regs0;
	xilinxmultiregimpl154_regs0 <= monroe_ionphoton_inj_o_sys50;
	xilinxmultiregimpl154_regs1 <= xilinxmultiregimpl154_regs0;
	xilinxmultiregimpl155_regs0 <= monroe_ionphoton_inj_o_sys51;
	xilinxmultiregimpl155_regs1 <= xilinxmultiregimpl155_regs0;
	xilinxmultiregimpl156_regs0 <= monroe_ionphoton_inj_o_sys52;
	xilinxmultiregimpl156_regs1 <= xilinxmultiregimpl156_regs0;
	xilinxmultiregimpl157_regs0 <= monroe_ionphoton_inj_o_sys53;
	xilinxmultiregimpl157_regs1 <= xilinxmultiregimpl157_regs0;
	xilinxmultiregimpl158_regs0 <= monroe_ionphoton_inj_o_sys54;
	xilinxmultiregimpl158_regs1 <= xilinxmultiregimpl158_regs0;
	xilinxmultiregimpl159_regs0 <= monroe_ionphoton_inj_o_sys55;
	xilinxmultiregimpl159_regs1 <= xilinxmultiregimpl159_regs0;
	xilinxmultiregimpl160_regs0 <= monroe_ionphoton_inj_o_sys56;
	xilinxmultiregimpl160_regs1 <= xilinxmultiregimpl160_regs0;
	xilinxmultiregimpl161_regs0 <= monroe_ionphoton_inj_o_sys57;
	xilinxmultiregimpl161_regs1 <= xilinxmultiregimpl161_regs0;
	xilinxmultiregimpl162_regs0 <= monroe_ionphoton_inj_o_sys58;
	xilinxmultiregimpl162_regs1 <= xilinxmultiregimpl162_regs0;
	xilinxmultiregimpl163_regs0 <= monroe_ionphoton_inj_o_sys59;
	xilinxmultiregimpl163_regs1 <= xilinxmultiregimpl163_regs0;
	xilinxmultiregimpl164_regs0 <= monroe_ionphoton_inj_o_sys60;
	xilinxmultiregimpl164_regs1 <= xilinxmultiregimpl164_regs0;
	xilinxmultiregimpl165_regs0 <= monroe_ionphoton_inj_o_sys61;
	xilinxmultiregimpl165_regs1 <= xilinxmultiregimpl165_regs0;
	xilinxmultiregimpl166_regs0 <= monroe_ionphoton_inj_o_sys62;
	xilinxmultiregimpl166_regs1 <= xilinxmultiregimpl166_regs0;
	xilinxmultiregimpl167_regs0 <= monroe_ionphoton_inj_o_sys63;
	xilinxmultiregimpl167_regs1 <= xilinxmultiregimpl167_regs0;
	xilinxmultiregimpl168_regs0 <= monroe_ionphoton_inj_o_sys64;
	xilinxmultiregimpl168_regs1 <= xilinxmultiregimpl168_regs0;
	xilinxmultiregimpl169_regs0 <= monroe_ionphoton_inj_o_sys65;
	xilinxmultiregimpl169_regs1 <= xilinxmultiregimpl169_regs0;
	xilinxmultiregimpl170_regs0 <= monroe_ionphoton_inj_o_sys66;
	xilinxmultiregimpl170_regs1 <= xilinxmultiregimpl170_regs0;
	xilinxmultiregimpl171_regs0 <= monroe_ionphoton_inj_o_sys67;
	xilinxmultiregimpl171_regs1 <= xilinxmultiregimpl171_regs0;
	xilinxmultiregimpl172_regs0 <= monroe_ionphoton_inj_o_sys68;
	xilinxmultiregimpl172_regs1 <= xilinxmultiregimpl172_regs0;
	xilinxmultiregimpl173_regs0 <= monroe_ionphoton_inj_o_sys69;
	xilinxmultiregimpl173_regs1 <= xilinxmultiregimpl173_regs0;
end

always @(posedge rio_phy_clk) begin
	if ((inout_8x0_inout_8x0_ointerface0_stb & (inout_8x0_inout_8x0_ointerface0_address == 1'd1))) begin
		inout_8x0_inout_8x0_oe_k <= inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (inout_8x0_inout_8x0_override_en) begin
		inout_8x0_serdes_oe <= inout_8x0_inout_8x0_override_oe;
	end else begin
		inout_8x0_serdes_oe <= inout_8x0_inout_8x0_oe_k;
	end
	inout_8x0_inout_8x0_i_d <= inout_8x0_serdes_i0[7];
	inout_8x0_inout_8x0_iinterface0_stb <= ((inout_8x0_inout_8x0_sample | (inout_8x0_inout_8x0_sensitivity[0] & (inout_8x0_serdes_i0[7] & (~inout_8x0_inout_8x0_i_d)))) | (inout_8x0_inout_8x0_sensitivity[1] & ((~inout_8x0_serdes_i0[7]) & inout_8x0_inout_8x0_i_d)));
	inout_8x0_inout_8x0_iinterface0_data <= inout_8x0_serdes_i0[7];
	inout_8x0_inout_8x0_iinterface0_fine_ts <= inout_8x0_inout_8x0_o;
	if ((inout_8x0_inout_8x0_ointerface0_stb & (inout_8x0_inout_8x0_ointerface0_address == 1'd0))) begin
		inout_8x0_inout_8x0_previous_data <= inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (inout_8x0_inout_8x0_override_en) begin
		inout_8x0_serdes_o0 <= {8{inout_8x0_inout_8x0_override_o}};
	end else begin
		if ((((inout_8x0_inout_8x0_ointerface0_stb & (inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & (~inout_8x0_inout_8x0_previous_data)) & inout_8x0_inout_8x0_ointerface0_data[0])) begin
			inout_8x0_serdes_o0 <= sync_f_t_array_muxed1;
		end else begin
			if ((((inout_8x0_inout_8x0_ointerface0_stb & (inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & inout_8x0_inout_8x0_previous_data) & (~inout_8x0_inout_8x0_ointerface0_data[0]))) begin
				inout_8x0_serdes_o0 <= sync_f_t_array_muxed2;
			end else begin
				inout_8x0_serdes_o0 <= {8{inout_8x0_inout_8x0_previous_data}};
			end
		end
	end
	if ((inout_8x1_inout_8x1_ointerface1_stb & (inout_8x1_inout_8x1_ointerface1_address == 1'd1))) begin
		inout_8x1_inout_8x1_oe_k <= inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (inout_8x1_inout_8x1_override_en) begin
		inout_8x1_serdes_oe <= inout_8x1_inout_8x1_override_oe;
	end else begin
		inout_8x1_serdes_oe <= inout_8x1_inout_8x1_oe_k;
	end
	inout_8x1_inout_8x1_i_d <= inout_8x1_serdes_i0[7];
	inout_8x1_inout_8x1_iinterface1_stb <= ((inout_8x1_inout_8x1_sample | (inout_8x1_inout_8x1_sensitivity[0] & (inout_8x1_serdes_i0[7] & (~inout_8x1_inout_8x1_i_d)))) | (inout_8x1_inout_8x1_sensitivity[1] & ((~inout_8x1_serdes_i0[7]) & inout_8x1_inout_8x1_i_d)));
	inout_8x1_inout_8x1_iinterface1_data <= inout_8x1_serdes_i0[7];
	inout_8x1_inout_8x1_iinterface1_fine_ts <= inout_8x1_inout_8x1_o;
	if ((inout_8x1_inout_8x1_ointerface1_stb & (inout_8x1_inout_8x1_ointerface1_address == 1'd0))) begin
		inout_8x1_inout_8x1_previous_data <= inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (inout_8x1_inout_8x1_override_en) begin
		inout_8x1_serdes_o0 <= {8{inout_8x1_inout_8x1_override_o}};
	end else begin
		if ((((inout_8x1_inout_8x1_ointerface1_stb & (inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & (~inout_8x1_inout_8x1_previous_data)) & inout_8x1_inout_8x1_ointerface1_data[0])) begin
			inout_8x1_serdes_o0 <= sync_f_t_array_muxed3;
		end else begin
			if ((((inout_8x1_inout_8x1_ointerface1_stb & (inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & inout_8x1_inout_8x1_previous_data) & (~inout_8x1_inout_8x1_ointerface1_data[0]))) begin
				inout_8x1_serdes_o0 <= sync_f_t_array_muxed4;
			end else begin
				inout_8x1_serdes_o0 <= {8{inout_8x1_inout_8x1_previous_data}};
			end
		end
	end
	if ((inout_8x2_inout_8x2_ointerface2_stb & (inout_8x2_inout_8x2_ointerface2_address == 1'd1))) begin
		inout_8x2_inout_8x2_oe_k <= inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (inout_8x2_inout_8x2_override_en) begin
		inout_8x2_serdes_oe <= inout_8x2_inout_8x2_override_oe;
	end else begin
		inout_8x2_serdes_oe <= inout_8x2_inout_8x2_oe_k;
	end
	inout_8x2_inout_8x2_i_d <= inout_8x2_serdes_i0[7];
	inout_8x2_inout_8x2_iinterface2_stb <= ((inout_8x2_inout_8x2_sample | (inout_8x2_inout_8x2_sensitivity[0] & (inout_8x2_serdes_i0[7] & (~inout_8x2_inout_8x2_i_d)))) | (inout_8x2_inout_8x2_sensitivity[1] & ((~inout_8x2_serdes_i0[7]) & inout_8x2_inout_8x2_i_d)));
	inout_8x2_inout_8x2_iinterface2_data <= inout_8x2_serdes_i0[7];
	inout_8x2_inout_8x2_iinterface2_fine_ts <= inout_8x2_inout_8x2_o;
	if ((inout_8x2_inout_8x2_ointerface2_stb & (inout_8x2_inout_8x2_ointerface2_address == 1'd0))) begin
		inout_8x2_inout_8x2_previous_data <= inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (inout_8x2_inout_8x2_override_en) begin
		inout_8x2_serdes_o0 <= {8{inout_8x2_inout_8x2_override_o}};
	end else begin
		if ((((inout_8x2_inout_8x2_ointerface2_stb & (inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & (~inout_8x2_inout_8x2_previous_data)) & inout_8x2_inout_8x2_ointerface2_data[0])) begin
			inout_8x2_serdes_o0 <= sync_f_t_array_muxed5;
		end else begin
			if ((((inout_8x2_inout_8x2_ointerface2_stb & (inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & inout_8x2_inout_8x2_previous_data) & (~inout_8x2_inout_8x2_ointerface2_data[0]))) begin
				inout_8x2_serdes_o0 <= sync_f_t_array_muxed6;
			end else begin
				inout_8x2_serdes_o0 <= {8{inout_8x2_inout_8x2_previous_data}};
			end
		end
	end
	if ((inout_8x3_inout_8x3_ointerface3_stb & (inout_8x3_inout_8x3_ointerface3_address == 1'd1))) begin
		inout_8x3_inout_8x3_oe_k <= inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (inout_8x3_inout_8x3_override_en) begin
		inout_8x3_serdes_oe <= inout_8x3_inout_8x3_override_oe;
	end else begin
		inout_8x3_serdes_oe <= inout_8x3_inout_8x3_oe_k;
	end
	inout_8x3_inout_8x3_i_d <= inout_8x3_serdes_i0[7];
	inout_8x3_inout_8x3_iinterface3_stb <= ((inout_8x3_inout_8x3_sample | (inout_8x3_inout_8x3_sensitivity[0] & (inout_8x3_serdes_i0[7] & (~inout_8x3_inout_8x3_i_d)))) | (inout_8x3_inout_8x3_sensitivity[1] & ((~inout_8x3_serdes_i0[7]) & inout_8x3_inout_8x3_i_d)));
	inout_8x3_inout_8x3_iinterface3_data <= inout_8x3_serdes_i0[7];
	inout_8x3_inout_8x3_iinterface3_fine_ts <= inout_8x3_inout_8x3_o;
	if ((inout_8x3_inout_8x3_ointerface3_stb & (inout_8x3_inout_8x3_ointerface3_address == 1'd0))) begin
		inout_8x3_inout_8x3_previous_data <= inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (inout_8x3_inout_8x3_override_en) begin
		inout_8x3_serdes_o0 <= {8{inout_8x3_inout_8x3_override_o}};
	end else begin
		if ((((inout_8x3_inout_8x3_ointerface3_stb & (inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & (~inout_8x3_inout_8x3_previous_data)) & inout_8x3_inout_8x3_ointerface3_data[0])) begin
			inout_8x3_serdes_o0 <= sync_f_t_array_muxed7;
		end else begin
			if ((((inout_8x3_inout_8x3_ointerface3_stb & (inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & inout_8x3_inout_8x3_previous_data) & (~inout_8x3_inout_8x3_ointerface3_data[0]))) begin
				inout_8x3_serdes_o0 <= sync_f_t_array_muxed8;
			end else begin
				inout_8x3_serdes_o0 <= {8{inout_8x3_inout_8x3_previous_data}};
			end
		end
	end
	if (output_8x0_stb) begin
		output_8x0_previous_data <= output_8x0_data;
	end
	if (output_8x0_override_en) begin
		output_8x0_o <= {8{output_8x0_override_o}};
	end else begin
		if (((output_8x0_stb & (~output_8x0_previous_data)) & output_8x0_data)) begin
			output_8x0_o <= sync_f_t_array_muxed9;
		end else begin
			if (((output_8x0_stb & output_8x0_previous_data) & (~output_8x0_data))) begin
				output_8x0_o <= sync_f_t_array_muxed10;
			end else begin
				output_8x0_o <= {8{output_8x0_previous_data}};
			end
		end
	end
	if (output_8x1_stb) begin
		output_8x1_previous_data <= output_8x1_data;
	end
	if (output_8x1_override_en) begin
		output_8x1_o <= {8{output_8x1_override_o}};
	end else begin
		if (((output_8x1_stb & (~output_8x1_previous_data)) & output_8x1_data)) begin
			output_8x1_o <= sync_f_t_array_muxed11;
		end else begin
			if (((output_8x1_stb & output_8x1_previous_data) & (~output_8x1_data))) begin
				output_8x1_o <= sync_f_t_array_muxed12;
			end else begin
				output_8x1_o <= {8{output_8x1_previous_data}};
			end
		end
	end
	if (output_8x2_stb) begin
		output_8x2_previous_data <= output_8x2_data;
	end
	if (output_8x2_override_en) begin
		output_8x2_o <= {8{output_8x2_override_o}};
	end else begin
		if (((output_8x2_stb & (~output_8x2_previous_data)) & output_8x2_data)) begin
			output_8x2_o <= sync_f_t_array_muxed13;
		end else begin
			if (((output_8x2_stb & output_8x2_previous_data) & (~output_8x2_data))) begin
				output_8x2_o <= sync_f_t_array_muxed14;
			end else begin
				output_8x2_o <= {8{output_8x2_previous_data}};
			end
		end
	end
	if (output_8x3_stb) begin
		output_8x3_previous_data <= output_8x3_data;
	end
	if (output_8x3_override_en) begin
		output_8x3_o <= {8{output_8x3_override_o}};
	end else begin
		if (((output_8x3_stb & (~output_8x3_previous_data)) & output_8x3_data)) begin
			output_8x3_o <= sync_f_t_array_muxed15;
		end else begin
			if (((output_8x3_stb & output_8x3_previous_data) & (~output_8x3_data))) begin
				output_8x3_o <= sync_f_t_array_muxed16;
			end else begin
				output_8x3_o <= {8{output_8x3_previous_data}};
			end
		end
	end
	if (output_8x4_stb) begin
		output_8x4_previous_data <= output_8x4_data;
	end
	if (output_8x4_override_en) begin
		output_8x4_o <= {8{output_8x4_override_o}};
	end else begin
		if (((output_8x4_stb & (~output_8x4_previous_data)) & output_8x4_data)) begin
			output_8x4_o <= sync_f_t_array_muxed17;
		end else begin
			if (((output_8x4_stb & output_8x4_previous_data) & (~output_8x4_data))) begin
				output_8x4_o <= sync_f_t_array_muxed18;
			end else begin
				output_8x4_o <= {8{output_8x4_previous_data}};
			end
		end
	end
	if (output_8x5_stb) begin
		output_8x5_previous_data <= output_8x5_data;
	end
	if (output_8x5_override_en) begin
		output_8x5_o <= {8{output_8x5_override_o}};
	end else begin
		if (((output_8x5_stb & (~output_8x5_previous_data)) & output_8x5_data)) begin
			output_8x5_o <= sync_f_t_array_muxed19;
		end else begin
			if (((output_8x5_stb & output_8x5_previous_data) & (~output_8x5_data))) begin
				output_8x5_o <= sync_f_t_array_muxed20;
			end else begin
				output_8x5_o <= {8{output_8x5_previous_data}};
			end
		end
	end
	if (output_8x6_stb) begin
		output_8x6_previous_data <= output_8x6_data;
	end
	if (output_8x6_override_en) begin
		output_8x6_o <= {8{output_8x6_override_o}};
	end else begin
		if (((output_8x6_stb & (~output_8x6_previous_data)) & output_8x6_data)) begin
			output_8x6_o <= sync_f_t_array_muxed21;
		end else begin
			if (((output_8x6_stb & output_8x6_previous_data) & (~output_8x6_data))) begin
				output_8x6_o <= sync_f_t_array_muxed22;
			end else begin
				output_8x6_o <= {8{output_8x6_previous_data}};
			end
		end
	end
	if (output_8x7_stb) begin
		output_8x7_previous_data <= output_8x7_data;
	end
	if (output_8x7_override_en) begin
		output_8x7_o <= {8{output_8x7_override_o}};
	end else begin
		if (((output_8x7_stb & (~output_8x7_previous_data)) & output_8x7_data)) begin
			output_8x7_o <= sync_f_t_array_muxed23;
		end else begin
			if (((output_8x7_stb & output_8x7_previous_data) & (~output_8x7_data))) begin
				output_8x7_o <= sync_f_t_array_muxed24;
			end else begin
				output_8x7_o <= {8{output_8x7_previous_data}};
			end
		end
	end
	if (output_8x8_stb) begin
		output_8x8_previous_data <= output_8x8_data;
	end
	if (output_8x8_override_en) begin
		output_8x8_o <= {8{output_8x8_override_o}};
	end else begin
		if (((output_8x8_stb & (~output_8x8_previous_data)) & output_8x8_data)) begin
			output_8x8_o <= sync_f_t_array_muxed25;
		end else begin
			if (((output_8x8_stb & output_8x8_previous_data) & (~output_8x8_data))) begin
				output_8x8_o <= sync_f_t_array_muxed26;
			end else begin
				output_8x8_o <= {8{output_8x8_previous_data}};
			end
		end
	end
	if (output_8x9_stb) begin
		output_8x9_previous_data <= output_8x9_data;
	end
	if (output_8x9_override_en) begin
		output_8x9_o <= {8{output_8x9_override_o}};
	end else begin
		if (((output_8x9_stb & (~output_8x9_previous_data)) & output_8x9_data)) begin
			output_8x9_o <= sync_f_t_array_muxed27;
		end else begin
			if (((output_8x9_stb & output_8x9_previous_data) & (~output_8x9_data))) begin
				output_8x9_o <= sync_f_t_array_muxed28;
			end else begin
				output_8x9_o <= {8{output_8x9_previous_data}};
			end
		end
	end
	if (output_8x10_stb) begin
		output_8x10_previous_data <= output_8x10_data;
	end
	if (output_8x10_override_en) begin
		output_8x10_o <= {8{output_8x10_override_o}};
	end else begin
		if (((output_8x10_stb & (~output_8x10_previous_data)) & output_8x10_data)) begin
			output_8x10_o <= sync_f_t_array_muxed29;
		end else begin
			if (((output_8x10_stb & output_8x10_previous_data) & (~output_8x10_data))) begin
				output_8x10_o <= sync_f_t_array_muxed30;
			end else begin
				output_8x10_o <= {8{output_8x10_previous_data}};
			end
		end
	end
	if (output_8x11_stb) begin
		output_8x11_previous_data <= output_8x11_data;
	end
	if (output_8x11_override_en) begin
		output_8x11_o <= {8{output_8x11_override_o}};
	end else begin
		if (((output_8x11_stb & (~output_8x11_previous_data)) & output_8x11_data)) begin
			output_8x11_o <= sync_f_t_array_muxed31;
		end else begin
			if (((output_8x11_stb & output_8x11_previous_data) & (~output_8x11_data))) begin
				output_8x11_o <= sync_f_t_array_muxed32;
			end else begin
				output_8x11_o <= {8{output_8x11_previous_data}};
			end
		end
	end
	if (spimaster0_iinterface0_stb) begin
		spimaster0_read <= 1'd0;
	end
	if ((spimaster0_ointerface0_stb & spimaster0_spimachine0_writable)) begin
		if (spimaster0_ointerface0_address) begin
			{spimaster0_config_cs, spimaster0_config_div, spimaster0_config_padding, spimaster0_config_length, spimaster0_config_half_duplex, spimaster0_config_lsb_first, spimaster0_config_clk_phase, spimaster0_config_clk_polarity, spimaster0_config_cs_polarity, spimaster0_config_input, spimaster0_config_end, spimaster0_config_offline} <= spimaster0_ointerface0_data;
		end else begin
			spimaster0_read <= spimaster0_config_input;
		end
	end
	if (spimaster0_interface_ce) begin
		spimaster0_interface_cs1 <= (({3{spimaster0_interface_cs_next}} & spimaster0_interface_cs0) ^ (~spimaster0_interface_cs_polarity));
		spimaster0_interface_clk <= (spimaster0_interface_clk_next ^ spimaster0_interface_clk_polarity);
	end
	if (spimaster0_interface_sample) begin
		spimaster0_interface_miso_reg <= spimaster0_interface_miso;
		spimaster0_interface_mosi_reg <= spimaster0_interface_mosi;
	end
	if (spimaster0_spimachine0_load1) begin
		spimaster0_spimachine0_n <= spimaster0_spimachine0_length;
		spimaster0_spimachine0_end1 <= spimaster0_spimachine0_end0;
	end
	if (spimaster0_spimachine0_shift) begin
		spimaster0_spimachine0_n <= (spimaster0_spimachine0_n - 1'd1);
	end
	if (spimaster0_spimachine0_shift) begin
		spimaster0_spimachine0_sr <= spimaster0_spimachine0_pdi;
		spimaster0_spimachine0_sdo <= (spimaster0_spimachine0_lsb_first ? spimaster0_spimachine0_pdi[0] : spimaster0_spimachine0_pdi[31]);
	end
	if (spimaster0_spimachine0_load1) begin
		spimaster0_spimachine0_sr <= spimaster0_spimachine0_pdo;
		spimaster0_spimachine0_sdo <= (spimaster0_spimachine0_lsb_first ? spimaster0_spimachine0_pdo[0] : spimaster0_spimachine0_pdo[31]);
	end
	if (spimaster0_spimachine0_count) begin
		if (spimaster0_spimachine0_cnt_done) begin
			if (spimaster0_spimachine0_do_extend) begin
				spimaster0_spimachine0_do_extend <= 1'd0;
			end else begin
				spimaster0_spimachine0_cnt <= spimaster0_spimachine0_div[7:1];
				spimaster0_spimachine0_do_extend <= (spimaster0_spimachine0_extend & spimaster0_spimachine0_div[0]);
			end
		end else begin
			spimaster0_spimachine0_cnt <= (spimaster0_spimachine0_cnt - 1'd1);
		end
	end
	spimaster0_state <= spimaster0_next_state;
	if (output_8x12_stb) begin
		output_8x12_previous_data <= output_8x12_data;
	end
	if (output_8x12_override_en) begin
		output_8x12_o <= {8{output_8x12_override_o}};
	end else begin
		if (((output_8x12_stb & (~output_8x12_previous_data)) & output_8x12_data)) begin
			output_8x12_o <= sync_f_t_array_muxed33;
		end else begin
			if (((output_8x12_stb & output_8x12_previous_data) & (~output_8x12_data))) begin
				output_8x12_o <= sync_f_t_array_muxed34;
			end else begin
				output_8x12_o <= {8{output_8x12_previous_data}};
			end
		end
	end
	if (output_8x13_stb) begin
		output_8x13_previous_data <= output_8x13_data;
	end
	if (output_8x13_override_en) begin
		output_8x13_o <= {8{output_8x13_override_o}};
	end else begin
		if (((output_8x13_stb & (~output_8x13_previous_data)) & output_8x13_data)) begin
			output_8x13_o <= sync_f_t_array_muxed35;
		end else begin
			if (((output_8x13_stb & output_8x13_previous_data) & (~output_8x13_data))) begin
				output_8x13_o <= sync_f_t_array_muxed36;
			end else begin
				output_8x13_o <= {8{output_8x13_previous_data}};
			end
		end
	end
	if (output_8x14_stb) begin
		output_8x14_previous_data <= output_8x14_data;
	end
	if (output_8x14_override_en) begin
		output_8x14_o <= {8{output_8x14_override_o}};
	end else begin
		if (((output_8x14_stb & (~output_8x14_previous_data)) & output_8x14_data)) begin
			output_8x14_o <= sync_f_t_array_muxed37;
		end else begin
			if (((output_8x14_stb & output_8x14_previous_data) & (~output_8x14_data))) begin
				output_8x14_o <= sync_f_t_array_muxed38;
			end else begin
				output_8x14_o <= {8{output_8x14_previous_data}};
			end
		end
	end
	if (output_8x15_stb) begin
		output_8x15_previous_data <= output_8x15_data;
	end
	if (output_8x15_override_en) begin
		output_8x15_o <= {8{output_8x15_override_o}};
	end else begin
		if (((output_8x15_stb & (~output_8x15_previous_data)) & output_8x15_data)) begin
			output_8x15_o <= sync_f_t_array_muxed39;
		end else begin
			if (((output_8x15_stb & output_8x15_previous_data) & (~output_8x15_data))) begin
				output_8x15_o <= sync_f_t_array_muxed40;
			end else begin
				output_8x15_o <= {8{output_8x15_previous_data}};
			end
		end
	end
	if (output_8x16_stb) begin
		output_8x16_previous_data <= output_8x16_data;
	end
	if (output_8x16_override_en) begin
		output_8x16_o <= {8{output_8x16_override_o}};
	end else begin
		if (((output_8x16_stb & (~output_8x16_previous_data)) & output_8x16_data)) begin
			output_8x16_o <= sync_f_t_array_muxed41;
		end else begin
			if (((output_8x16_stb & output_8x16_previous_data) & (~output_8x16_data))) begin
				output_8x16_o <= sync_f_t_array_muxed42;
			end else begin
				output_8x16_o <= {8{output_8x16_previous_data}};
			end
		end
	end
	if (spimaster1_iinterface1_stb) begin
		spimaster1_read <= 1'd0;
	end
	if ((spimaster1_ointerface1_stb & spimaster1_spimachine1_writable)) begin
		if (spimaster1_ointerface1_address) begin
			{spimaster1_config_cs, spimaster1_config_div, spimaster1_config_padding, spimaster1_config_length, spimaster1_config_half_duplex, spimaster1_config_lsb_first, spimaster1_config_clk_phase, spimaster1_config_clk_polarity, spimaster1_config_cs_polarity, spimaster1_config_input, spimaster1_config_end, spimaster1_config_offline} <= spimaster1_ointerface1_data;
		end else begin
			spimaster1_read <= spimaster1_config_input;
		end
	end
	if (spimaster1_interface_ce) begin
		spimaster1_interface_cs1 <= (({3{spimaster1_interface_cs_next}} & spimaster1_interface_cs0) ^ (~spimaster1_interface_cs_polarity));
		spimaster1_interface_clk <= (spimaster1_interface_clk_next ^ spimaster1_interface_clk_polarity);
	end
	if (spimaster1_interface_sample) begin
		spimaster1_interface_miso_reg <= spimaster1_interface_miso;
		spimaster1_interface_mosi_reg <= spimaster1_interface_mosi;
	end
	if (spimaster1_spimachine1_load1) begin
		spimaster1_spimachine1_n <= spimaster1_spimachine1_length;
		spimaster1_spimachine1_end1 <= spimaster1_spimachine1_end0;
	end
	if (spimaster1_spimachine1_shift) begin
		spimaster1_spimachine1_n <= (spimaster1_spimachine1_n - 1'd1);
	end
	if (spimaster1_spimachine1_shift) begin
		spimaster1_spimachine1_sr <= spimaster1_spimachine1_pdi;
		spimaster1_spimachine1_sdo <= (spimaster1_spimachine1_lsb_first ? spimaster1_spimachine1_pdi[0] : spimaster1_spimachine1_pdi[31]);
	end
	if (spimaster1_spimachine1_load1) begin
		spimaster1_spimachine1_sr <= spimaster1_spimachine1_pdo;
		spimaster1_spimachine1_sdo <= (spimaster1_spimachine1_lsb_first ? spimaster1_spimachine1_pdo[0] : spimaster1_spimachine1_pdo[31]);
	end
	if (spimaster1_spimachine1_count) begin
		if (spimaster1_spimachine1_cnt_done) begin
			if (spimaster1_spimachine1_do_extend) begin
				spimaster1_spimachine1_do_extend <= 1'd0;
			end else begin
				spimaster1_spimachine1_cnt <= spimaster1_spimachine1_div[7:1];
				spimaster1_spimachine1_do_extend <= (spimaster1_spimachine1_extend & spimaster1_spimachine1_div[0]);
			end
		end else begin
			spimaster1_spimachine1_cnt <= (spimaster1_spimachine1_cnt - 1'd1);
		end
	end
	spimaster1_state <= spimaster1_next_state;
	if (output_8x17_stb) begin
		output_8x17_previous_data <= output_8x17_data;
	end
	if (output_8x17_override_en) begin
		output_8x17_o <= {8{output_8x17_override_o}};
	end else begin
		if (((output_8x17_stb & (~output_8x17_previous_data)) & output_8x17_data)) begin
			output_8x17_o <= sync_f_t_array_muxed43;
		end else begin
			if (((output_8x17_stb & output_8x17_previous_data) & (~output_8x17_data))) begin
				output_8x17_o <= sync_f_t_array_muxed44;
			end else begin
				output_8x17_o <= {8{output_8x17_previous_data}};
			end
		end
	end
	if (output_8x18_stb) begin
		output_8x18_previous_data <= output_8x18_data;
	end
	if (output_8x18_override_en) begin
		output_8x18_o <= {8{output_8x18_override_o}};
	end else begin
		if (((output_8x18_stb & (~output_8x18_previous_data)) & output_8x18_data)) begin
			output_8x18_o <= sync_f_t_array_muxed45;
		end else begin
			if (((output_8x18_stb & output_8x18_previous_data) & (~output_8x18_data))) begin
				output_8x18_o <= sync_f_t_array_muxed46;
			end else begin
				output_8x18_o <= {8{output_8x18_previous_data}};
			end
		end
	end
	if (output_8x19_stb) begin
		output_8x19_previous_data <= output_8x19_data;
	end
	if (output_8x19_override_en) begin
		output_8x19_o <= {8{output_8x19_override_o}};
	end else begin
		if (((output_8x19_stb & (~output_8x19_previous_data)) & output_8x19_data)) begin
			output_8x19_o <= sync_f_t_array_muxed47;
		end else begin
			if (((output_8x19_stb & output_8x19_previous_data) & (~output_8x19_data))) begin
				output_8x19_o <= sync_f_t_array_muxed48;
			end else begin
				output_8x19_o <= {8{output_8x19_previous_data}};
			end
		end
	end
	if (output_8x20_stb) begin
		output_8x20_previous_data <= output_8x20_data;
	end
	if (output_8x20_override_en) begin
		output_8x20_o <= {8{output_8x20_override_o}};
	end else begin
		if (((output_8x20_stb & (~output_8x20_previous_data)) & output_8x20_data)) begin
			output_8x20_o <= sync_f_t_array_muxed49;
		end else begin
			if (((output_8x20_stb & output_8x20_previous_data) & (~output_8x20_data))) begin
				output_8x20_o <= sync_f_t_array_muxed50;
			end else begin
				output_8x20_o <= {8{output_8x20_previous_data}};
			end
		end
	end
	if (output_8x21_stb) begin
		output_8x21_previous_data <= output_8x21_data;
	end
	if (output_8x21_override_en) begin
		output_8x21_o <= {8{output_8x21_override_o}};
	end else begin
		if (((output_8x21_stb & (~output_8x21_previous_data)) & output_8x21_data)) begin
			output_8x21_o <= sync_f_t_array_muxed51;
		end else begin
			if (((output_8x21_stb & output_8x21_previous_data) & (~output_8x21_data))) begin
				output_8x21_o <= sync_f_t_array_muxed52;
			end else begin
				output_8x21_o <= {8{output_8x21_previous_data}};
			end
		end
	end
	if (spimaster2_iinterface2_stb) begin
		spimaster2_read <= 1'd0;
	end
	if ((spimaster2_ointerface2_stb & spimaster2_spimachine2_writable)) begin
		if (spimaster2_ointerface2_address) begin
			{spimaster2_config_cs, spimaster2_config_div, spimaster2_config_padding, spimaster2_config_length, spimaster2_config_half_duplex, spimaster2_config_lsb_first, spimaster2_config_clk_phase, spimaster2_config_clk_polarity, spimaster2_config_cs_polarity, spimaster2_config_input, spimaster2_config_end, spimaster2_config_offline} <= spimaster2_ointerface2_data;
		end else begin
			spimaster2_read <= spimaster2_config_input;
		end
	end
	if (spimaster2_interface_ce) begin
		spimaster2_interface_cs1 <= (({3{spimaster2_interface_cs_next}} & spimaster2_interface_cs0) ^ (~spimaster2_interface_cs_polarity));
		spimaster2_interface_clk <= (spimaster2_interface_clk_next ^ spimaster2_interface_clk_polarity);
	end
	if (spimaster2_interface_sample) begin
		spimaster2_interface_miso_reg <= spimaster2_interface_miso;
		spimaster2_interface_mosi_reg <= spimaster2_interface_mosi;
	end
	if (spimaster2_spimachine2_load1) begin
		spimaster2_spimachine2_n <= spimaster2_spimachine2_length;
		spimaster2_spimachine2_end1 <= spimaster2_spimachine2_end0;
	end
	if (spimaster2_spimachine2_shift) begin
		spimaster2_spimachine2_n <= (spimaster2_spimachine2_n - 1'd1);
	end
	if (spimaster2_spimachine2_shift) begin
		spimaster2_spimachine2_sr <= spimaster2_spimachine2_pdi;
		spimaster2_spimachine2_sdo <= (spimaster2_spimachine2_lsb_first ? spimaster2_spimachine2_pdi[0] : spimaster2_spimachine2_pdi[31]);
	end
	if (spimaster2_spimachine2_load1) begin
		spimaster2_spimachine2_sr <= spimaster2_spimachine2_pdo;
		spimaster2_spimachine2_sdo <= (spimaster2_spimachine2_lsb_first ? spimaster2_spimachine2_pdo[0] : spimaster2_spimachine2_pdo[31]);
	end
	if (spimaster2_spimachine2_count) begin
		if (spimaster2_spimachine2_cnt_done) begin
			if (spimaster2_spimachine2_do_extend) begin
				spimaster2_spimachine2_do_extend <= 1'd0;
			end else begin
				spimaster2_spimachine2_cnt <= spimaster2_spimachine2_div[7:1];
				spimaster2_spimachine2_do_extend <= (spimaster2_spimachine2_extend & spimaster2_spimachine2_div[0]);
			end
		end else begin
			spimaster2_spimachine2_cnt <= (spimaster2_spimachine2_cnt - 1'd1);
		end
	end
	spimaster2_state <= spimaster2_next_state;
	if (output_8x22_stb) begin
		output_8x22_previous_data <= output_8x22_data;
	end
	if (output_8x22_override_en) begin
		output_8x22_o <= {8{output_8x22_override_o}};
	end else begin
		if (((output_8x22_stb & (~output_8x22_previous_data)) & output_8x22_data)) begin
			output_8x22_o <= sync_f_t_array_muxed53;
		end else begin
			if (((output_8x22_stb & output_8x22_previous_data) & (~output_8x22_data))) begin
				output_8x22_o <= sync_f_t_array_muxed54;
			end else begin
				output_8x22_o <= {8{output_8x22_previous_data}};
			end
		end
	end
	if (output_8x23_stb) begin
		output_8x23_previous_data <= output_8x23_data;
	end
	if (output_8x23_override_en) begin
		output_8x23_o <= {8{output_8x23_override_o}};
	end else begin
		if (((output_8x23_stb & (~output_8x23_previous_data)) & output_8x23_data)) begin
			output_8x23_o <= sync_f_t_array_muxed55;
		end else begin
			if (((output_8x23_stb & output_8x23_previous_data) & (~output_8x23_data))) begin
				output_8x23_o <= sync_f_t_array_muxed56;
			end else begin
				output_8x23_o <= {8{output_8x23_previous_data}};
			end
		end
	end
	if (output_8x24_stb) begin
		output_8x24_previous_data <= output_8x24_data;
	end
	if (output_8x24_override_en) begin
		output_8x24_o <= {8{output_8x24_override_o}};
	end else begin
		if (((output_8x24_stb & (~output_8x24_previous_data)) & output_8x24_data)) begin
			output_8x24_o <= sync_f_t_array_muxed57;
		end else begin
			if (((output_8x24_stb & output_8x24_previous_data) & (~output_8x24_data))) begin
				output_8x24_o <= sync_f_t_array_muxed58;
			end else begin
				output_8x24_o <= {8{output_8x24_previous_data}};
			end
		end
	end
	if (output_8x25_stb) begin
		output_8x25_previous_data <= output_8x25_data;
	end
	if (output_8x25_override_en) begin
		output_8x25_o <= {8{output_8x25_override_o}};
	end else begin
		if (((output_8x25_stb & (~output_8x25_previous_data)) & output_8x25_data)) begin
			output_8x25_o <= sync_f_t_array_muxed59;
		end else begin
			if (((output_8x25_stb & output_8x25_previous_data) & (~output_8x25_data))) begin
				output_8x25_o <= sync_f_t_array_muxed60;
			end else begin
				output_8x25_o <= {8{output_8x25_previous_data}};
			end
		end
	end
	if (output_8x26_stb) begin
		output_8x26_previous_data <= output_8x26_data;
	end
	if (output_8x26_override_en) begin
		output_8x26_o <= {8{output_8x26_override_o}};
	end else begin
		if (((output_8x26_stb & (~output_8x26_previous_data)) & output_8x26_data)) begin
			output_8x26_o <= sync_f_t_array_muxed61;
		end else begin
			if (((output_8x26_stb & output_8x26_previous_data) & (~output_8x26_data))) begin
				output_8x26_o <= sync_f_t_array_muxed62;
			end else begin
				output_8x26_o <= {8{output_8x26_previous_data}};
			end
		end
	end
	if (output0_stb) begin
		output0_pad_k <= output0_data;
	end
	if (output0_override_en) begin
		output0_pad_o <= output0_override_o;
	end else begin
		output0_pad_o <= output0_pad_k;
	end
	if (output1_stb) begin
		output1_pad_k <= output1_data;
	end
	if (output1_override_en) begin
		output1_pad_o <= output1_override_o;
	end else begin
		output1_pad_o <= output1_pad_k;
	end
	if (rio_phy_rst) begin
		inout_8x0_serdes_o0 <= 8'd0;
		inout_8x0_serdes_oe <= 1'd0;
		inout_8x0_inout_8x0_iinterface0_stb <= 1'd0;
		inout_8x0_inout_8x0_previous_data <= 1'd0;
		inout_8x0_inout_8x0_oe_k <= 1'd0;
		inout_8x0_inout_8x0_i_d <= 1'd0;
		inout_8x1_serdes_o0 <= 8'd0;
		inout_8x1_serdes_oe <= 1'd0;
		inout_8x1_inout_8x1_iinterface1_stb <= 1'd0;
		inout_8x1_inout_8x1_previous_data <= 1'd0;
		inout_8x1_inout_8x1_oe_k <= 1'd0;
		inout_8x1_inout_8x1_i_d <= 1'd0;
		inout_8x2_serdes_o0 <= 8'd0;
		inout_8x2_serdes_oe <= 1'd0;
		inout_8x2_inout_8x2_iinterface2_stb <= 1'd0;
		inout_8x2_inout_8x2_previous_data <= 1'd0;
		inout_8x2_inout_8x2_oe_k <= 1'd0;
		inout_8x2_inout_8x2_i_d <= 1'd0;
		inout_8x3_serdes_o0 <= 8'd0;
		inout_8x3_serdes_oe <= 1'd0;
		inout_8x3_inout_8x3_iinterface3_stb <= 1'd0;
		inout_8x3_inout_8x3_previous_data <= 1'd0;
		inout_8x3_inout_8x3_oe_k <= 1'd0;
		inout_8x3_inout_8x3_i_d <= 1'd0;
		output_8x0_o <= 8'd0;
		output_8x0_previous_data <= 1'd0;
		output_8x1_o <= 8'd0;
		output_8x1_previous_data <= 1'd0;
		output_8x2_o <= 8'd0;
		output_8x2_previous_data <= 1'd0;
		output_8x3_o <= 8'd0;
		output_8x3_previous_data <= 1'd0;
		output_8x4_o <= 8'd0;
		output_8x4_previous_data <= 1'd0;
		output_8x5_o <= 8'd0;
		output_8x5_previous_data <= 1'd0;
		output_8x6_o <= 8'd0;
		output_8x6_previous_data <= 1'd0;
		output_8x7_o <= 8'd0;
		output_8x7_previous_data <= 1'd0;
		output_8x8_o <= 8'd0;
		output_8x8_previous_data <= 1'd0;
		output_8x9_o <= 8'd0;
		output_8x9_previous_data <= 1'd0;
		output_8x10_o <= 8'd0;
		output_8x10_previous_data <= 1'd0;
		output_8x11_o <= 8'd0;
		output_8x11_previous_data <= 1'd0;
		spimaster0_interface_cs1 <= 3'd7;
		spimaster0_interface_clk <= 1'd0;
		spimaster0_spimachine0_cnt <= 7'd0;
		spimaster0_spimachine0_do_extend <= 1'd0;
		spimaster0_config_offline <= 1'd1;
		spimaster0_config_end <= 1'd1;
		spimaster0_config_input <= 1'd0;
		spimaster0_config_cs_polarity <= 1'd0;
		spimaster0_config_clk_polarity <= 1'd0;
		spimaster0_config_clk_phase <= 1'd0;
		spimaster0_config_lsb_first <= 1'd0;
		spimaster0_config_half_duplex <= 1'd0;
		spimaster0_config_length <= 5'd0;
		spimaster0_config_padding <= 3'd0;
		spimaster0_config_div <= 8'd0;
		spimaster0_config_cs <= 8'd0;
		spimaster0_read <= 1'd0;
		output_8x12_o <= 8'd0;
		output_8x12_previous_data <= 1'd0;
		output_8x13_o <= 8'd0;
		output_8x13_previous_data <= 1'd0;
		output_8x14_o <= 8'd0;
		output_8x14_previous_data <= 1'd0;
		output_8x15_o <= 8'd0;
		output_8x15_previous_data <= 1'd0;
		output_8x16_o <= 8'd0;
		output_8x16_previous_data <= 1'd0;
		spimaster1_interface_cs1 <= 3'd7;
		spimaster1_interface_clk <= 1'd0;
		spimaster1_spimachine1_cnt <= 7'd0;
		spimaster1_spimachine1_do_extend <= 1'd0;
		spimaster1_config_offline <= 1'd1;
		spimaster1_config_end <= 1'd1;
		spimaster1_config_input <= 1'd0;
		spimaster1_config_cs_polarity <= 1'd0;
		spimaster1_config_clk_polarity <= 1'd0;
		spimaster1_config_clk_phase <= 1'd0;
		spimaster1_config_lsb_first <= 1'd0;
		spimaster1_config_half_duplex <= 1'd0;
		spimaster1_config_length <= 5'd0;
		spimaster1_config_padding <= 3'd0;
		spimaster1_config_div <= 8'd0;
		spimaster1_config_cs <= 8'd0;
		spimaster1_read <= 1'd0;
		output_8x17_o <= 8'd0;
		output_8x17_previous_data <= 1'd0;
		output_8x18_o <= 8'd0;
		output_8x18_previous_data <= 1'd0;
		output_8x19_o <= 8'd0;
		output_8x19_previous_data <= 1'd0;
		output_8x20_o <= 8'd0;
		output_8x20_previous_data <= 1'd0;
		output_8x21_o <= 8'd0;
		output_8x21_previous_data <= 1'd0;
		spimaster2_interface_cs1 <= 3'd7;
		spimaster2_interface_clk <= 1'd0;
		spimaster2_spimachine2_cnt <= 7'd0;
		spimaster2_spimachine2_do_extend <= 1'd0;
		spimaster2_config_offline <= 1'd1;
		spimaster2_config_end <= 1'd1;
		spimaster2_config_input <= 1'd0;
		spimaster2_config_cs_polarity <= 1'd0;
		spimaster2_config_clk_polarity <= 1'd0;
		spimaster2_config_clk_phase <= 1'd0;
		spimaster2_config_lsb_first <= 1'd0;
		spimaster2_config_half_duplex <= 1'd0;
		spimaster2_config_length <= 5'd0;
		spimaster2_config_padding <= 3'd0;
		spimaster2_config_div <= 8'd0;
		spimaster2_config_cs <= 8'd0;
		spimaster2_read <= 1'd0;
		output_8x22_o <= 8'd0;
		output_8x22_previous_data <= 1'd0;
		output_8x23_o <= 8'd0;
		output_8x23_previous_data <= 1'd0;
		output_8x24_o <= 8'd0;
		output_8x24_previous_data <= 1'd0;
		output_8x25_o <= 8'd0;
		output_8x25_previous_data <= 1'd0;
		output_8x26_o <= 8'd0;
		output_8x26_previous_data <= 1'd0;
		output0_pad_k <= 1'd0;
		output1_pad_k <= 1'd0;
		spimaster0_state <= 3'd0;
		spimaster1_state <= 3'd0;
		spimaster2_state <= 3'd0;
	end
end

always @(posedge rsys_clk) begin
	monroe_ionphoton_rtio_core_outputs_lanedistributor_min_minus_timestamp <= (monroe_ionphoton_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp);
	monroe_ionphoton_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp <= (sync_rhs_array_muxed3 - monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp);
	monroe_ionphoton_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp <= (sync_rhs_array_muxed4 - monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp);
	monroe_ionphoton_rtio_core_outputs_lanedistributor_last_minus_timestamp <= (monroe_ionphoton_rtio_core_outputs_lanedistributor_last_coarse_timestamp - monroe_ionphoton_rtio_core_outputs_lanedistributor_coarse_timestamp);
	monroe_ionphoton_rtio_core_outputs_lanedistributor_quash <= 1'd0;
	if ((monroe_ionphoton_rtio_core_cri_chan_sel[15:0] == 6'd36)) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_quash <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane <= monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		sync_t_lhs_array_muxed = monroe_ionphoton_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		case (monroe_ionphoton_rtio_core_outputs_lanedistributor_use_lanen)
			1'd0: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= sync_t_lhs_array_muxed;
			end
			1'd1: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= sync_t_lhs_array_muxed;
			end
			2'd2: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= sync_t_lhs_array_muxed;
			end
			2'd3: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= sync_t_lhs_array_muxed;
			end
			3'd4: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= sync_t_lhs_array_muxed;
			end
			3'd5: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= sync_t_lhs_array_muxed;
			end
			3'd6: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= sync_t_lhs_array_muxed;
			end
			default: begin
				monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= sync_t_lhs_array_muxed;
			end
		endcase
		monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn <= (monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn + 1'd1);
	end
	if ((monroe_ionphoton_rtio_core_cri_cmd == 1'd1)) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_outputs_lanedistributor_do_underflow) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd1;
	end
	monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error <= monroe_ionphoton_rtio_core_outputs_lanedistributor_do_sequence_error;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error_channel <= monroe_ionphoton_rtio_core_cri_chan_sel[15:0];
	monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable_r <= monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable;
	if (((~monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable_r) & monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable)) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_force_laneB <= 1'd1;
	end
	if (monroe_ionphoton_rtio_core_outputs_lanedistributor_do_write) begin
		monroe_ionphoton_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
	end
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
	monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
	if ((monroe_ionphoton_rtio_core_inputs_selected0 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow0 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer0_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow0 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected1 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow1 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer1_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow1 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected2 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow2 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer2_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow2 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected3 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow3 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer3_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow3 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected4 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow4 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer4_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow4 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected5 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow5 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer5_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow5 <= 1'd1;
	end
	if ((monroe_ionphoton_rtio_core_inputs_selected6 & monroe_ionphoton_rtio_core_inputs_i_ack)) begin
		monroe_ionphoton_rtio_core_inputs_overflow6 <= 1'd0;
	end
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer6_o) begin
		monroe_ionphoton_rtio_core_inputs_overflow6 <= 1'd1;
	end
	monroe_ionphoton_rtio_core_inputs_i_ack <= 1'd0;
	if (monroe_ionphoton_rtio_core_inputs_i_ack) begin
		monroe_ionphoton_rtio_core_cri_i_status <= {1'd0, monroe_ionphoton_rtio_core_inputs_i_status_raw[1], (~monroe_ionphoton_rtio_core_inputs_i_status_raw[0])};
		monroe_ionphoton_rtio_core_cri_i_data <= sync_t_rhs_array_muxed1;
		monroe_ionphoton_rtio_core_cri_i_timestamp <= sync_t_rhs_array_muxed2;
	end
	if (((monroe_ionphoton_rtio_tsc_full_ts_sys >= monroe_ionphoton_rtio_core_inputs_input_timeout) | (monroe_ionphoton_rtio_core_inputs_i_status_raw != 1'd0))) begin
		if (monroe_ionphoton_rtio_core_inputs_input_pending) begin
			monroe_ionphoton_rtio_core_inputs_i_ack <= 1'd1;
		end
		monroe_ionphoton_rtio_core_inputs_input_pending <= 1'd0;
	end
	if ((monroe_ionphoton_rtio_core_cri_cmd == 2'd2)) begin
		monroe_ionphoton_rtio_core_inputs_input_timeout <= monroe_ionphoton_rtio_core_cri_i_timeout;
		monroe_ionphoton_rtio_core_inputs_input_pending <= 1'd1;
		monroe_ionphoton_rtio_core_cri_i_status <= 3'd4;
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
	monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
	monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o_r <= monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_i) begin
		monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o_r <= monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_i) begin
		monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_o_collision_sync_ps_ack_toggle_i);
	end
	monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o_r <= monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_o;
	if (monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_i) begin
		monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_i <= (~monroe_ionphoton_rtio_core_o_busy_sync_ps_ack_toggle_i);
	end
	if (rsys_rst) begin
		monroe_ionphoton_rtio_core_cri_i_status <= 4'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane <= 3'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= 61'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_seqn <= 12'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_quash <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_current_lane_writable_r <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= 8'd0;
		monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= 8'd0;
		monroe_ionphoton_rtio_core_inputs_i_ack <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_overflow0 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_overflow1 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_overflow2 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= 7'd0;
		monroe_ionphoton_rtio_core_inputs_overflow3 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_overflow4 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_overflow5 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= 3'd0;
		monroe_ionphoton_rtio_core_inputs_overflow6 <= 1'd0;
		monroe_ionphoton_rtio_core_inputs_input_pending <= 1'd0;
	end
	xilinxmultiregimpl18_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_graycounter1_q;
	xilinxmultiregimpl18_regs1 <= xilinxmultiregimpl18_regs0;
	xilinxmultiregimpl20_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_graycounter3_q;
	xilinxmultiregimpl20_regs1 <= xilinxmultiregimpl20_regs0;
	xilinxmultiregimpl22_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_graycounter5_q;
	xilinxmultiregimpl22_regs1 <= xilinxmultiregimpl22_regs0;
	xilinxmultiregimpl24_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_graycounter7_q;
	xilinxmultiregimpl24_regs1 <= xilinxmultiregimpl24_regs0;
	xilinxmultiregimpl26_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_graycounter9_q;
	xilinxmultiregimpl26_regs1 <= xilinxmultiregimpl26_regs0;
	xilinxmultiregimpl28_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_graycounter11_q;
	xilinxmultiregimpl28_regs1 <= xilinxmultiregimpl28_regs0;
	xilinxmultiregimpl30_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_graycounter13_q;
	xilinxmultiregimpl30_regs1 <= xilinxmultiregimpl30_regs0;
	xilinxmultiregimpl32_regs0 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_graycounter15_q;
	xilinxmultiregimpl32_regs1 <= xilinxmultiregimpl32_regs0;
	xilinxmultiregimpl33_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_graycounter0_q;
	xilinxmultiregimpl33_regs1 <= xilinxmultiregimpl33_regs0;
	xilinxmultiregimpl35_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer0_ps_toggle_i;
	xilinxmultiregimpl35_regs1 <= xilinxmultiregimpl35_regs0;
	xilinxmultiregimpl37_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_graycounter2_q;
	xilinxmultiregimpl37_regs1 <= xilinxmultiregimpl37_regs0;
	xilinxmultiregimpl39_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer1_ps_toggle_i;
	xilinxmultiregimpl39_regs1 <= xilinxmultiregimpl39_regs0;
	xilinxmultiregimpl41_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_graycounter4_q;
	xilinxmultiregimpl41_regs1 <= xilinxmultiregimpl41_regs0;
	xilinxmultiregimpl43_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer2_ps_toggle_i;
	xilinxmultiregimpl43_regs1 <= xilinxmultiregimpl43_regs0;
	xilinxmultiregimpl45_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_graycounter6_q;
	xilinxmultiregimpl45_regs1 <= xilinxmultiregimpl45_regs0;
	xilinxmultiregimpl47_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer3_ps_toggle_i;
	xilinxmultiregimpl47_regs1 <= xilinxmultiregimpl47_regs0;
	xilinxmultiregimpl49_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_graycounter8_q;
	xilinxmultiregimpl49_regs1 <= xilinxmultiregimpl49_regs0;
	xilinxmultiregimpl51_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer4_ps_toggle_i;
	xilinxmultiregimpl51_regs1 <= xilinxmultiregimpl51_regs0;
	xilinxmultiregimpl53_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_graycounter10_q;
	xilinxmultiregimpl53_regs1 <= xilinxmultiregimpl53_regs0;
	xilinxmultiregimpl55_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer5_ps_toggle_i;
	xilinxmultiregimpl55_regs1 <= xilinxmultiregimpl55_regs0;
	xilinxmultiregimpl57_regs0 <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_graycounter12_q;
	xilinxmultiregimpl57_regs1 <= xilinxmultiregimpl57_regs0;
	xilinxmultiregimpl59_regs0 <= monroe_ionphoton_rtio_core_inputs_blindtransfer6_ps_toggle_i;
	xilinxmultiregimpl59_regs1 <= xilinxmultiregimpl59_regs0;
	xilinxmultiregimpl61_regs0 <= monroe_ionphoton_rtio_core_o_collision_sync_ps_toggle_i;
	xilinxmultiregimpl61_regs1 <= xilinxmultiregimpl61_regs0;
	xilinxmultiregimpl63_regs0 <= monroe_ionphoton_rtio_core_o_collision_sync_bxfer_data;
	xilinxmultiregimpl63_regs1 <= xilinxmultiregimpl63_regs0;
	xilinxmultiregimpl64_regs0 <= monroe_ionphoton_rtio_core_o_busy_sync_ps_toggle_i;
	xilinxmultiregimpl64_regs1 <= xilinxmultiregimpl64_regs0;
	xilinxmultiregimpl66_regs0 <= monroe_ionphoton_rtio_core_o_busy_sync_bxfer_data;
	xilinxmultiregimpl66_regs1 <= xilinxmultiregimpl66_regs0;
end

always @(posedge rtio_clk) begin
	if (monroe_ionphoton_rtio_tsc_load) begin
		monroe_ionphoton_rtio_tsc_coarse_ts <= monroe_ionphoton_rtio_tsc_load_value;
	end else begin
		monroe_ionphoton_rtio_tsc_coarse_ts <= (monroe_ionphoton_rtio_tsc_coarse_ts + 1'd1);
	end
	monroe_ionphoton_rtio_tsc_value_gray_rtio <= (monroe_ionphoton_rtio_tsc_i ^ monroe_ionphoton_rtio_tsc_i[60:1]);
	if (rtio_rst) begin
		monroe_ionphoton_rtio_tsc_coarse_ts <= 61'd0;
	end
end

always @(posedge sys_clk) begin
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_adr[29:10] == 1'd0))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error <= 1'd1;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_adr[29:10] == monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_stb) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_w;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_adr;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_r;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter == 1'd1)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_we;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter == 2'd2)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_ack <= 1'd1;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter == 2'd3)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_ack <= 1'd0;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter != 1'd0)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter + 1'd1);
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_stb)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter <= 1'd1;
		end
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_stb & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy)) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_payload_data;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_txen & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount + 1'd1);
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy <= 1'd0;
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack <= 1'd1;
				end else begin
					serial_tx <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg[0];
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg <= {1'd0, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy) begin
		{monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_txen, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_tx} <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_tx + monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage);
	end else begin
		{monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_txen, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_stb <= 1'd0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx;
	if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy)) begin
		if (((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_r)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy <= 1'd1;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_rxen) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount + 1'd1);
			if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount == 1'd0)) begin
				if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx) begin
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount == 4'd9)) begin
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy <= 1'd0;
					if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx) begin
						monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_payload_data <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_reg;
						monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_stb <= 1'd1;
					end
				end else begin
					monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_reg <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy) begin
		{monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_rxen, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_rx} <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_rx + monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage);
	end else begin
		{monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_rxen, monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_clear) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_pending <= 1'd0;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_old_trigger <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_trigger;
	if (((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_trigger) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_old_trigger)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_pending <= 1'd1;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_clear) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_pending <= 1'd0;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_old_trigger <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_trigger;
	if (((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_trigger) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_old_trigger)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_pending <= 1'd1;
	end
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_replace))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce + 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_do_read) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_consume <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_consume + 1'd1);
	end
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_replace))) begin
		if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_do_read)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_do_read) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_replace))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce + 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_do_read) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_consume <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_consume + 1'd1);
	end
	if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_replace))) begin
		if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_do_read)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_do_read) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level - 1'd1);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage) begin
		if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value == 1'd0)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage;
		end else begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value - 1'd1);
		end
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_clear) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_pending <= 1'd0;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_old_trigger <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_trigger;
	if (((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_trigger) & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_old_trigger)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_pending <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en0 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_en;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en0;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en2 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en1;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en3 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en2;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en3;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_valid <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en[2:0], monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_en};
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dqs <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe;
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata_valid) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p0_rddata;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata_valid) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p1_rddata;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata_valid) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p2_rddata;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata_valid) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_inti_p3_rddata;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce0) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset0) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce1) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset1) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce2) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset2) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce3) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset3) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce4) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset4) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce5) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset5) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce6) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset6) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_ce7) begin
		if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_open) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle <= 1'd0;
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row0;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_reset7) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row1 <= 15'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_wait) begin
		if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_done)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count - 1'd1);
		end
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count <= 3'd4;
	end
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_wait) begin
		if ((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_done)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count - 1'd1);
		end
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count <= 10'd886;
	end
	minicon_state <= minicon_next_state;
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_adr_offset_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_cpulevel_sdram_if_arbitrated_adr[1:0];
	fullmemorywe_state <= fullmemorywe_next_state;
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 == 1'd0)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_clk <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dqi <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i0;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 == 1'd1)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_clk <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr[29:0], monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dqi};
	end else begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 + 1'd1);
	end
	if ((((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_stb) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 == 1'd1)) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 1'd0))) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dq_oe <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_cs_n <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr[31:16] <= 16'd61423;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 5'd16)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr[31:8] <= {monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_adr, {2{1'd0}}};
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 6'd40)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dq_oe <= 1'd0;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 7'd82)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_ack <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_cs_n <= 1'd1;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 7'd83)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_ack <= 1'd0;
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 7'd85)) begin
	end
	if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter == 7'd85)) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter != 1'd0)) begin
			monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter <= (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter + 1'd1);
		end else begin
			if (((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_cyc & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_stb) & (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 == 1'd1))) begin
				monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter <= 1'd1;
			end
		end
	end
	monroe_ionphoton_monroe_ionphoton_tx_mmcm_reset <= (~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_lock);
	if (monroe_ionphoton_monroe_ionphoton_rx_reset) begin
		monroe_ionphoton_monroe_ionphoton_cdr_locked <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_cdr_lock_counter <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_cdr_lock_counter != 13'd4531)) begin
			monroe_ionphoton_monroe_ionphoton_cdr_lock_counter <= (monroe_ionphoton_monroe_ionphoton_cdr_lock_counter + 1'd1);
		end else begin
			monroe_ionphoton_monroe_ionphoton_cdr_locked <= 1'd1;
		end
	end
	monroe_ionphoton_monroe_ionphoton_rx_mmcm_reset <= (~monroe_ionphoton_monroe_ionphoton_cdr_locked);
	monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset0 <= monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset1;
	monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset0 <= monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset1;
	monroe_ionphoton_monroe_ionphoton_tx_init_tick <= 1'd0;
	if ((monroe_ionphoton_monroe_ionphoton_tx_init_timer == 6'd57)) begin
		monroe_ionphoton_monroe_ionphoton_tx_init_tick <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_tx_init_timer <= 1'd0;
	end else begin
		monroe_ionphoton_monroe_ionphoton_tx_init_timer <= (monroe_ionphoton_monroe_ionphoton_tx_init_timer + 1'd1);
	end
	a7_1000basex_gtptxinit_state <= a7_1000basex_gtptxinit_next_state;
	monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset0 <= monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset1;
	monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done_r <= monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done1;
	a7_1000basex_gtprxinit_state <= a7_1000basex_gtprxinit_next_state;
	if (monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value_ce) begin
		monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue <= monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue_gtprxinit_next_value;
	end
	monroe_ionphoton_monroe_ionphoton_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_toggle_o;
	if (monroe_ionphoton_monroe_ionphoton_ps_preamble_error_o) begin
		monroe_ionphoton_monroe_ionphoton_preamble_errors_status <= (monroe_ionphoton_monroe_ionphoton_preamble_errors_status + 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_ps_crc_error_o) begin
		monroe_ionphoton_monroe_ionphoton_crc_errors_status <= (monroe_ionphoton_monroe_ionphoton_crc_errors_status + 1'd1);
	end
	monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_o;
	monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o_r <= monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_o;
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next_binary;
	monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_next;
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_binary <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next_binary;
	monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_next;
	if (monroe_ionphoton_monroe_ionphoton_writer_counter_reset) begin
		monroe_ionphoton_monroe_ionphoton_writer_counter <= 1'd0;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_writer_counter_ce) begin
			monroe_ionphoton_monroe_ionphoton_writer_counter <= (monroe_ionphoton_monroe_ionphoton_writer_counter + monroe_ionphoton_monroe_ionphoton_writer_increment);
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_writer_slot_ce) begin
		monroe_ionphoton_monroe_ionphoton_writer_slot <= (monroe_ionphoton_monroe_ionphoton_writer_slot + 1'd1);
	end
	if (((monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_writer_fifo_replace))) begin
		monroe_ionphoton_monroe_ionphoton_writer_fifo_produce <= (monroe_ionphoton_monroe_ionphoton_writer_fifo_produce + 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_writer_fifo_do_read) begin
		monroe_ionphoton_monroe_ionphoton_writer_fifo_consume <= (monroe_ionphoton_monroe_ionphoton_writer_fifo_consume + 1'd1);
	end
	if (((monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_writer_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_writer_fifo_replace))) begin
		if ((~monroe_ionphoton_monroe_ionphoton_writer_fifo_do_read)) begin
			monroe_ionphoton_monroe_ionphoton_writer_fifo_level <= (monroe_ionphoton_monroe_ionphoton_writer_fifo_level + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_writer_fifo_do_read) begin
			monroe_ionphoton_monroe_ionphoton_writer_fifo_level <= (monroe_ionphoton_monroe_ionphoton_writer_fifo_level - 1'd1);
		end
	end
	liteethmacsramwriter_state <= liteethmacsramwriter_next_state;
	if (monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value_ce) begin
		monroe_ionphoton_monroe_ionphoton_writer_errors_status <= monroe_ionphoton_monroe_ionphoton_writer_errors_status_next_value;
	end
	if (monroe_ionphoton_monroe_ionphoton_reader_counter_reset) begin
		monroe_ionphoton_monroe_ionphoton_reader_counter <= 1'd0;
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_reader_counter_ce) begin
			monroe_ionphoton_monroe_ionphoton_reader_counter <= (monroe_ionphoton_monroe_ionphoton_reader_counter + 3'd4);
		end
	end
	monroe_ionphoton_monroe_ionphoton_reader_last_d <= monroe_ionphoton_monroe_ionphoton_reader_last;
	if (monroe_ionphoton_monroe_ionphoton_reader_done_clear) begin
		monroe_ionphoton_monroe_ionphoton_reader_done_pending <= 1'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_reader_done_trigger) begin
		monroe_ionphoton_monroe_ionphoton_reader_done_pending <= 1'd1;
	end
	if (((monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_reader_fifo_replace))) begin
		monroe_ionphoton_monroe_ionphoton_reader_fifo_produce <= (monroe_ionphoton_monroe_ionphoton_reader_fifo_produce + 1'd1);
	end
	if (monroe_ionphoton_monroe_ionphoton_reader_fifo_do_read) begin
		monroe_ionphoton_monroe_ionphoton_reader_fifo_consume <= (monroe_ionphoton_monroe_ionphoton_reader_fifo_consume + 1'd1);
	end
	if (((monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_we & monroe_ionphoton_monroe_ionphoton_reader_fifo_syncfifo_writable) & (~monroe_ionphoton_monroe_ionphoton_reader_fifo_replace))) begin
		if ((~monroe_ionphoton_monroe_ionphoton_reader_fifo_do_read)) begin
			monroe_ionphoton_monroe_ionphoton_reader_fifo_level <= (monroe_ionphoton_monroe_ionphoton_reader_fifo_level + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_monroe_ionphoton_reader_fifo_do_read) begin
			monroe_ionphoton_monroe_ionphoton_reader_fifo_level <= (monroe_ionphoton_monroe_ionphoton_reader_fifo_level - 1'd1);
		end
	end
	liteethmacsramreader_state <= liteethmacsramreader_next_state;
	monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc0 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb0) & (~monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0))) begin
		monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc0 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb0) & (~monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0))) begin
		monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc0 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb0) & (~monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0))) begin
		monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc0 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb0) & (~monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0))) begin
		monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram0_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram0_bus_stb1) & (~monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1))) begin
		monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram1_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram1_bus_stb1) & (~monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1))) begin
		monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram2_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram2_bus_stb1) & (~monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1))) begin
		monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1 <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_sram3_bus_cyc1 & monroe_ionphoton_monroe_ionphoton_sram3_bus_stb1) & (~monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1))) begin
		monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1 <= 1'd1;
	end
	monroe_ionphoton_monroe_ionphoton_slave_sel_r <= monroe_ionphoton_monroe_ionphoton_slave_sel;
	case (grant)
		1'd0: begin
			if ((~request[0])) begin
				if (request[1]) begin
					grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~request[1])) begin
				if (request[0]) begin
					grant <= 1'd0;
				end
			end
		end
	endcase
	slave_sel_r <= slave_sel;
	monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_r <= sync_rhs_array_muxed5;
	monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_mailbox_i1_cyc & monroe_ionphoton_monroe_ionphoton_mailbox_i1_stb) & (~monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack))) begin
		monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack <= 1'd1;
		if (monroe_ionphoton_monroe_ionphoton_mailbox_i1_we) begin
			sync_t_t_array_muxed0 = monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_w;
			case (monroe_ionphoton_monroe_ionphoton_mailbox_i1_adr[1:0])
				1'd0: begin
					monroe_ionphoton_monroe_ionphoton_mailbox0 <= sync_t_t_array_muxed0;
				end
				1'd1: begin
					monroe_ionphoton_monroe_ionphoton_mailbox1 <= sync_t_t_array_muxed0;
				end
				default: begin
					monroe_ionphoton_monroe_ionphoton_mailbox2 <= sync_t_t_array_muxed0;
				end
			endcase
		end
	end
	monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_r <= sync_rhs_array_muxed6;
	monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack <= 1'd0;
	if (((monroe_ionphoton_monroe_ionphoton_mailbox_i2_cyc & monroe_ionphoton_monroe_ionphoton_mailbox_i2_stb) & (~monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack))) begin
		monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack <= 1'd1;
		if (monroe_ionphoton_monroe_ionphoton_mailbox_i2_we) begin
			sync_t_t_array_muxed1 = monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_w;
			case (monroe_ionphoton_monroe_ionphoton_mailbox_i2_adr[1:0])
				1'd0: begin
					monroe_ionphoton_monroe_ionphoton_mailbox0 <= sync_t_t_array_muxed1;
				end
				1'd1: begin
					monroe_ionphoton_monroe_ionphoton_mailbox1 <= sync_t_t_array_muxed1;
				end
				default: begin
					monroe_ionphoton_monroe_ionphoton_mailbox2 <= sync_t_t_array_muxed1;
				end
			endcase
		end
	end
	monroe_ionphoton_rtio_tsc_o <= monroe_ionphoton_rtio_tsc_value_sys;
	monroe_ionphoton_rtio_core_cmd_reset <= monroe_ionphoton_rtio_core_reset_re;
	monroe_ionphoton_rtio_core_cmd_reset_phy <= monroe_ionphoton_rtio_core_reset_phy_re;
	monroe_ionphoton_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= (monroe_ionphoton_rtio_tsc_coarse_ts_sys + 5'd16);
	if (monroe_ionphoton_rtio_core_async_error_re) begin
		if (monroe_ionphoton_rtio_core_async_error_r[0]) begin
			monroe_ionphoton_rtio_core_o_collision <= 1'd0;
		end
		if (monroe_ionphoton_rtio_core_async_error_r[1]) begin
			monroe_ionphoton_rtio_core_o_busy <= 1'd0;
		end
		if (monroe_ionphoton_rtio_core_async_error_r[2]) begin
			monroe_ionphoton_rtio_core_o_sequence_error <= 1'd0;
		end
	end
	if (monroe_ionphoton_rtio_core_o_collision_sync_o) begin
		monroe_ionphoton_rtio_core_o_collision <= 1'd1;
		if ((~monroe_ionphoton_rtio_core_o_collision)) begin
			monroe_ionphoton_rtio_core_collision_channel_status <= monroe_ionphoton_rtio_core_o_collision_sync_data_o;
		end
	end
	if (monroe_ionphoton_rtio_core_o_busy_sync_o) begin
		monroe_ionphoton_rtio_core_o_busy <= 1'd1;
		if ((~monroe_ionphoton_rtio_core_o_busy)) begin
			monroe_ionphoton_rtio_core_busy_channel_status <= monroe_ionphoton_rtio_core_o_busy_sync_data_o;
		end
	end
	if (monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error) begin
		monroe_ionphoton_rtio_core_o_sequence_error <= 1'd1;
		if ((~monroe_ionphoton_rtio_core_o_sequence_error)) begin
			monroe_ionphoton_rtio_core_sequence_error_channel_status <= monroe_ionphoton_rtio_core_outputs_lanedistributor_sequence_error_channel;
		end
	end
	if (monroe_ionphoton_rtio_now_hi_re) begin
		monroe_ionphoton_rtio_now_hi_backing <= monroe_ionphoton_rtio_now_hi_r;
	end
	if (monroe_ionphoton_rtio_now_lo_re) begin
		monroe_ionphoton_rtio_now <= {monroe_ionphoton_rtio_now_hi_backing, monroe_ionphoton_rtio_now_lo_r};
	end
	if (monroe_ionphoton_rtio_counter_update_re) begin
		monroe_ionphoton_rtio_counter_status <= monroe_ionphoton_rtio_tsc_full_ts_sys;
	end
	case (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_adr[4:0])
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_target0_w;
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_rtio_now_hi_w;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_rtio_now_lo_w;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_w;
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_w;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_w;
		end
		3'd6: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_w;
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_w;
		end
		4'd8: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_w;
		end
		4'd9: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_w;
		end
		4'd10: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_w;
		end
		4'd11: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_w;
		end
		4'd12: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_w;
		end
		4'd13: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_w;
		end
		4'd14: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_w;
		end
		4'd15: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_w;
		end
		5'd16: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_w;
		end
		5'd17: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_w;
		end
		5'd18: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_w;
		end
		5'd19: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_status_w;
		end
		5'd20: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_w;
		end
		5'd21: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_w;
		end
		5'd22: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_data_w;
		end
		5'd23: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp1_w;
		end
		5'd24: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timestamp0_w;
		end
		5'd25: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_status_w;
		end
		5'd26: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_rtio_i_overflow_reset_w;
		end
		5'd27: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_counter1_w;
		end
		5'd28: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank0_counter0_w;
		end
		5'd29: begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= monroe_ionphoton_rtio_counter_update_w;
		end
	endcase
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack) begin
		monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_csrbank0_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank0_bus_stb)) begin
			monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack <= 1'd1;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_target0_re) begin
		monroe_ionphoton_rtio_target_storage_full[31:0] <= monroe_ionphoton_monroe_ionphoton_csrbank0_target0_r;
	end
	monroe_ionphoton_rtio_target_re <= monroe_ionphoton_monroe_ionphoton_csrbank0_target0_re;
	if (monroe_ionphoton_rtio_o_data_we) begin
		monroe_ionphoton_rtio_o_data_storage_full <= (monroe_ionphoton_rtio_o_data_dat_w <<< 1'd0);
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[511:480] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data15_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[479:448] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data14_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[447:416] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data13_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[415:384] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data12_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[383:352] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data11_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[351:320] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data10_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[319:288] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data9_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[287:256] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data8_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[255:224] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data7_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[223:192] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data6_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[191:160] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data5_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[159:128] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data4_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[127:96] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data3_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[95:64] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data2_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[63:32] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data1_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_re) begin
		monroe_ionphoton_rtio_o_data_storage_full[31:0] <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_r;
	end
	monroe_ionphoton_rtio_o_data_re <= monroe_ionphoton_monroe_ionphoton_csrbank0_o_data0_re;
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_re) begin
		monroe_ionphoton_rtio_i_timeout_storage_full[63:32] <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout1_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_re) begin
		monroe_ionphoton_rtio_i_timeout_storage_full[31:0] <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_r;
	end
	monroe_ionphoton_rtio_i_timeout_re <= monroe_ionphoton_monroe_ionphoton_csrbank0_i_timeout0_re;
	case (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_adr[3:0])
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_dma_enable_enable_w;
		end
		1'd1: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_w;
		end
		2'd2: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_w;
		end
		2'd3: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_w;
		end
		3'd4: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_w;
		end
		3'd5: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_dma_cri_master_error_w;
		end
		3'd6: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_error_channel_w;
		end
		3'd7: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp1_w;
		end
		4'd8: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_error_timestamp0_w;
		end
		4'd9: begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank1_error_address_w;
		end
	endcase
	if (monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack) begin
		monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_csrbank1_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank1_bus_stb)) begin
			monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack <= 1'd1;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_re) begin
		monroe_ionphoton_dma_dma_storage_full[33:32] <= monroe_ionphoton_monroe_ionphoton_csrbank1_base_address1_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_re) begin
		monroe_ionphoton_dma_dma_storage_full[31:0] <= monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_r;
	end
	monroe_ionphoton_dma_dma_re <= monroe_ionphoton_monroe_ionphoton_csrbank1_base_address0_re;
	if (monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_re) begin
		monroe_ionphoton_dma_time_offset_storage_full[63:32] <= monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset1_r;
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_re) begin
		monroe_ionphoton_dma_time_offset_storage_full[31:0] <= monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_r;
	end
	monroe_ionphoton_dma_time_offset_re <= monroe_ionphoton_monroe_ionphoton_csrbank1_time_offset0_re;
	monroe_ionphoton_cri_con_selected <= monroe_ionphoton_cri_con_shared_chan_sel[23:16];
	case (monroe_ionphoton_monroe_ionphoton_csrbank2_bus_adr[0])
		1'd0: begin
			monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_w;
		end
	endcase
	if (monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack) begin
		monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack <= 1'd0;
	end else begin
		if ((monroe_ionphoton_monroe_ionphoton_csrbank2_bus_cyc & monroe_ionphoton_monroe_ionphoton_csrbank2_bus_stb)) begin
			monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack <= 1'd1;
		end
	end
	if (monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_re) begin
		monroe_ionphoton_cri_con_storage_full[1:0] <= monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_r;
	end
	monroe_ionphoton_cri_con_re <= monroe_ionphoton_monroe_ionphoton_csrbank2_selected0_re;
	if (monroe_ionphoton_mon_value_update_re) begin
		monroe_ionphoton_mon_status <= sync_t_rhs_array_muxed3;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd0)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys0 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd0)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys1 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd0)) & (monroe_ionphoton_inj_override_sel_storage == 2'd2))) begin
		monroe_ionphoton_inj_o_sys2 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd1)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys3 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd1)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys4 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 1'd1)) & (monroe_ionphoton_inj_override_sel_storage == 2'd2))) begin
		monroe_ionphoton_inj_o_sys5 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd2)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys6 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd2)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys7 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd2)) & (monroe_ionphoton_inj_override_sel_storage == 2'd2))) begin
		monroe_ionphoton_inj_o_sys8 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd3)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys9 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd3)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys10 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 2'd3)) & (monroe_ionphoton_inj_override_sel_storage == 2'd2))) begin
		monroe_ionphoton_inj_o_sys11 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd4)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys12 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd4)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys13 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd5)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys14 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd5)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys15 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd6)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys16 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd6)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys17 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd7)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys18 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 3'd7)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys19 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd8)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys20 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd8)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys21 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd9)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys22 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd9)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys23 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd10)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys24 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd10)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys25 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd11)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys26 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd11)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys27 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd12)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys28 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd12)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys29 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd13)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys30 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd13)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys31 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd14)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys32 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd14)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys33 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd15)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys34 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 4'd15)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys35 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd17)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys36 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd17)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys37 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd18)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys38 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd18)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys39 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd19)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys40 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd19)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys41 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd20)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys42 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd20)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys43 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd21)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys44 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd21)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys45 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd23)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys46 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd23)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys47 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd24)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys48 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd24)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys49 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd25)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys50 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd25)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys51 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd26)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys52 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd26)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys53 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd27)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys54 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd27)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys55 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd29)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys56 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd29)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys57 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd30)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys58 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd30)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys59 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd31)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys60 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 5'd31)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys61 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd32)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys62 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd32)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys63 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd33)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys64 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd33)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys65 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd34)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys66 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd34)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys67 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd35)) & (monroe_ionphoton_inj_override_sel_storage == 1'd0))) begin
		monroe_ionphoton_inj_o_sys68 <= monroe_ionphoton_inj_value_r;
	end
	if (((monroe_ionphoton_inj_value_re & (monroe_ionphoton_inj_chan_sel_storage == 6'd35)) & (monroe_ionphoton_inj_override_sel_storage == 1'd1))) begin
		monroe_ionphoton_inj_o_sys69 <= monroe_ionphoton_inj_value_r;
	end
	monroe_ionphoton_rtio_analyzer_enable_r <= monroe_ionphoton_rtio_analyzer_enable_storage;
	if ((monroe_ionphoton_rtio_analyzer_enable_storage & (~monroe_ionphoton_rtio_analyzer_enable_r))) begin
		monroe_ionphoton_rtio_analyzer_busy_status <= 1'd1;
	end
	if (((monroe_ionphoton_rtio_analyzer_dma_sink_stb & monroe_ionphoton_rtio_analyzer_dma_sink_ack) & monroe_ionphoton_rtio_analyzer_dma_sink_eop)) begin
		monroe_ionphoton_rtio_analyzer_busy_status <= 1'd0;
	end
	monroe_ionphoton_rtio_analyzer_message_encoder_read_wait_event_r <= monroe_ionphoton_rtio_core_cri_i_status[2];
	monroe_ionphoton_rtio_analyzer_message_encoder_just_written <= (monroe_ionphoton_rtio_core_cri_cmd == 1'd1);
	monroe_ionphoton_rtio_analyzer_message_encoder_enable_r <= monroe_ionphoton_rtio_analyzer_enable_storage;
	if (((~monroe_ionphoton_rtio_analyzer_enable_storage) & monroe_ionphoton_rtio_analyzer_message_encoder_enable_r)) begin
		monroe_ionphoton_rtio_analyzer_message_encoder_stopping <= 1'd1;
	end
	if ((~monroe_ionphoton_rtio_analyzer_message_encoder_stopping)) begin
		if (monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data <= {monroe_ionphoton_rtio_analyzer_message_encoder_exception_padding1, monroe_ionphoton_rtio_analyzer_message_encoder_exception_exception_type, monroe_ionphoton_rtio_analyzer_message_encoder_exception_rtio_counter, monroe_ionphoton_rtio_analyzer_message_encoder_exception_padding0, monroe_ionphoton_rtio_analyzer_message_encoder_exception_channel, monroe_ionphoton_rtio_analyzer_message_encoder_exception_message_type};
		end else begin
			monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data <= {monroe_ionphoton_rtio_analyzer_message_encoder_input_output_data, monroe_ionphoton_rtio_analyzer_message_encoder_input_output_address_padding, monroe_ionphoton_rtio_analyzer_message_encoder_input_output_rtio_counter, monroe_ionphoton_rtio_analyzer_message_encoder_input_output_timestamp, monroe_ionphoton_rtio_analyzer_message_encoder_input_output_channel, monroe_ionphoton_rtio_analyzer_message_encoder_input_output_message_type};
		end
		monroe_ionphoton_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_source_stb <= (monroe_ionphoton_rtio_analyzer_enable_storage & (monroe_ionphoton_rtio_analyzer_message_encoder_input_output_stb | monroe_ionphoton_rtio_analyzer_message_encoder_exception_stb));
		if (monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_re) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_status <= 1'd0;
		end
		if ((monroe_ionphoton_rtio_analyzer_message_encoder_source_stb & (~monroe_ionphoton_rtio_analyzer_message_encoder_source_ack))) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_status <= 1'd1;
		end
	end else begin
		monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data <= {monroe_ionphoton_rtio_analyzer_message_encoder_stopped_padding1, monroe_ionphoton_rtio_analyzer_message_encoder_stopped_rtio_counter, monroe_ionphoton_rtio_analyzer_message_encoder_stopped_padding0, monroe_ionphoton_rtio_analyzer_message_encoder_stopped_message_type};
		monroe_ionphoton_rtio_analyzer_message_encoder_source_eop <= 1'd1;
		monroe_ionphoton_rtio_analyzer_message_encoder_source_stb <= 1'd1;
		if (monroe_ionphoton_rtio_analyzer_message_encoder_source_ack) begin
			monroe_ionphoton_rtio_analyzer_message_encoder_stopping <= 1'd0;
		end
	end
	if (monroe_ionphoton_rtio_analyzer_fifo_syncfifo_re) begin
		monroe_ionphoton_rtio_analyzer_fifo_readable <= 1'd1;
	end else begin
		if (monroe_ionphoton_rtio_analyzer_fifo_re) begin
			monroe_ionphoton_rtio_analyzer_fifo_readable <= 1'd0;
		end
	end
	if (((monroe_ionphoton_rtio_analyzer_fifo_syncfifo_we & monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable) & (~monroe_ionphoton_rtio_analyzer_fifo_replace))) begin
		monroe_ionphoton_rtio_analyzer_fifo_produce <= (monroe_ionphoton_rtio_analyzer_fifo_produce + 1'd1);
	end
	if (monroe_ionphoton_rtio_analyzer_fifo_do_read) begin
		monroe_ionphoton_rtio_analyzer_fifo_consume <= (monroe_ionphoton_rtio_analyzer_fifo_consume + 1'd1);
	end
	if (((monroe_ionphoton_rtio_analyzer_fifo_syncfifo_we & monroe_ionphoton_rtio_analyzer_fifo_syncfifo_writable) & (~monroe_ionphoton_rtio_analyzer_fifo_replace))) begin
		if ((~monroe_ionphoton_rtio_analyzer_fifo_do_read)) begin
			monroe_ionphoton_rtio_analyzer_fifo_level0 <= (monroe_ionphoton_rtio_analyzer_fifo_level0 + 1'd1);
		end
	end else begin
		if (monroe_ionphoton_rtio_analyzer_fifo_do_read) begin
			monroe_ionphoton_rtio_analyzer_fifo_level0 <= (monroe_ionphoton_rtio_analyzer_fifo_level0 - 1'd1);
		end
	end
	if ((monroe_ionphoton_rtio_analyzer_converter_source_stb & monroe_ionphoton_rtio_analyzer_converter_source_ack)) begin
		if (monroe_ionphoton_rtio_analyzer_converter_last) begin
			monroe_ionphoton_rtio_analyzer_converter_mux <= 1'd0;
		end else begin
			monroe_ionphoton_rtio_analyzer_converter_mux <= (monroe_ionphoton_rtio_analyzer_converter_mux + 1'd1);
		end
	end
	if (monroe_ionphoton_rtio_analyzer_dma_reset_re) begin
		monroe_ionphoton_monroe_ionphoton_interface1_bus_adr <= monroe_ionphoton_rtio_analyzer_dma_base_address_storage;
	end
	if (monroe_ionphoton_monroe_ionphoton_interface1_bus_ack) begin
		if ((monroe_ionphoton_monroe_ionphoton_interface1_bus_adr == monroe_ionphoton_rtio_analyzer_dma_last_address_storage)) begin
			monroe_ionphoton_monroe_ionphoton_interface1_bus_adr <= monroe_ionphoton_rtio_analyzer_dma_base_address_storage;
		end else begin
			monroe_ionphoton_monroe_ionphoton_interface1_bus_adr <= (monroe_ionphoton_monroe_ionphoton_interface1_bus_adr + 1'd1);
		end
	end
	if (monroe_ionphoton_rtio_analyzer_dma_reset_re) begin
		monroe_ionphoton_rtio_analyzer_dma_message_count <= 1'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_interface1_bus_ack) begin
		monroe_ionphoton_rtio_analyzer_dma_message_count <= (monroe_ionphoton_rtio_analyzer_dma_message_count + monroe_ionphoton_rtio_analyzer_dma_sink_payload_valid_token_count);
	end
	case (sdram_cpulevel_arbiter_grant)
		1'd0: begin
			if ((~sdram_cpulevel_arbiter_request[0])) begin
				if (sdram_cpulevel_arbiter_request[1]) begin
					sdram_cpulevel_arbiter_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~sdram_cpulevel_arbiter_request[1])) begin
				if (sdram_cpulevel_arbiter_request[0]) begin
					sdram_cpulevel_arbiter_grant <= 1'd0;
				end
			end
		end
	endcase
	case (sdram_native_arbiter_grant)
		1'd0: begin
			if ((~sdram_native_arbiter_request[0])) begin
				if (sdram_native_arbiter_request[1]) begin
					sdram_native_arbiter_grant <= 1'd1;
				end else begin
					if (sdram_native_arbiter_request[2]) begin
						sdram_native_arbiter_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~sdram_native_arbiter_request[1])) begin
				if (sdram_native_arbiter_request[2]) begin
					sdram_native_arbiter_grant <= 2'd2;
				end else begin
					if (sdram_native_arbiter_request[0]) begin
						sdram_native_arbiter_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~sdram_native_arbiter_request[2])) begin
				if (sdram_native_arbiter_request[0]) begin
					sdram_native_arbiter_grant <= 1'd0;
				end else begin
					if (sdram_native_arbiter_request[1]) begin
						sdram_native_arbiter_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	case (monroe_ionphoton_grant)
		1'd0: begin
			if ((~monroe_ionphoton_request[0])) begin
				if (monroe_ionphoton_request[1]) begin
					monroe_ionphoton_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~monroe_ionphoton_request[1])) begin
				if (monroe_ionphoton_request[0]) begin
					monroe_ionphoton_grant <= 1'd0;
				end
			end
		end
	endcase
	monroe_ionphoton_slave_sel_r <= monroe_ionphoton_slave_sel;
	monroe_ionphoton_interface0_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank0_sel) begin
		case (monroe_ionphoton_interface0_bank_bus_adr[1:0])
			1'd0: begin
				monroe_ionphoton_interface0_bank_bus_dat_r <= monroe_ionphoton_csrbank0_dly_sel0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface0_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_w;
			end
			2'd2: begin
				monroe_ionphoton_interface0_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_w;
			end
			2'd3: begin
				monroe_ionphoton_interface0_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank0_dly_sel0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage_full[1:0] <= monroe_ionphoton_csrbank0_dly_sel0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_re <= monroe_ionphoton_csrbank0_dly_sel0_re;
	monroe_ionphoton_interface1_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank1_sel) begin
		case (monroe_ionphoton_interface1_bank_bus_adr[5:0])
			1'd0: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_control0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_command0_w;
			end
			2'd2: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_address1_w;
			end
			3'd4: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_address0_w;
			end
			3'd5: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_baddress0_w;
			end
			3'd6: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_wrdata3_w;
			end
			3'd7: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_wrdata2_w;
			end
			4'd8: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_wrdata1_w;
			end
			4'd9: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_wrdata0_w;
			end
			4'd10: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_rddata3_w;
			end
			4'd11: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_rddata2_w;
			end
			4'd12: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_rddata1_w;
			end
			4'd13: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi0_rddata0_w;
			end
			4'd14: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_command0_w;
			end
			4'd15: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_address1_w;
			end
			5'd17: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_address0_w;
			end
			5'd18: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_baddress0_w;
			end
			5'd19: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_wrdata3_w;
			end
			5'd20: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_wrdata2_w;
			end
			5'd21: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_wrdata1_w;
			end
			5'd22: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_wrdata0_w;
			end
			5'd23: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_rddata3_w;
			end
			5'd24: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_rddata2_w;
			end
			5'd25: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_rddata1_w;
			end
			5'd26: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi1_rddata0_w;
			end
			5'd27: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_command0_w;
			end
			5'd28: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_address1_w;
			end
			5'd30: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_address0_w;
			end
			5'd31: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_baddress0_w;
			end
			6'd32: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_wrdata3_w;
			end
			6'd33: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_wrdata2_w;
			end
			6'd34: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_wrdata1_w;
			end
			6'd35: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_wrdata0_w;
			end
			6'd36: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_rddata3_w;
			end
			6'd37: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_rddata2_w;
			end
			6'd38: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_rddata1_w;
			end
			6'd39: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi2_rddata0_w;
			end
			6'd40: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_command0_w;
			end
			6'd41: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_address1_w;
			end
			6'd43: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_address0_w;
			end
			6'd44: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_baddress0_w;
			end
			6'd45: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_wrdata3_w;
			end
			6'd46: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_wrdata2_w;
			end
			6'd47: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_wrdata1_w;
			end
			6'd48: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_wrdata0_w;
			end
			6'd49: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_rddata3_w;
			end
			6'd50: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_rddata2_w;
			end
			6'd51: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_rddata1_w;
			end
			6'd52: begin
				monroe_ionphoton_interface1_bank_bus_dat_r <= monroe_ionphoton_csrbank1_pi3_rddata0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank1_control0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage_full[3:0] <= monroe_ionphoton_csrbank1_control0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_re <= monroe_ionphoton_csrbank1_control0_re;
	if (monroe_ionphoton_csrbank1_pi0_command0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage_full[5:0] <= monroe_ionphoton_csrbank1_pi0_command0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_re <= monroe_ionphoton_csrbank1_pi0_command0_re;
	if (monroe_ionphoton_csrbank1_pi0_address1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full[14:8] <= monroe_ionphoton_csrbank1_pi0_address1_r;
	end
	if (monroe_ionphoton_csrbank1_pi0_address0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi0_address0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_re <= monroe_ionphoton_csrbank1_pi0_address0_re;
	if (monroe_ionphoton_csrbank1_pi0_baddress0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage_full[2:0] <= monroe_ionphoton_csrbank1_pi0_baddress0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_re <= monroe_ionphoton_csrbank1_pi0_baddress0_re;
	if (monroe_ionphoton_csrbank1_pi0_wrdata3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[31:24] <= monroe_ionphoton_csrbank1_pi0_wrdata3_r;
	end
	if (monroe_ionphoton_csrbank1_pi0_wrdata2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[23:16] <= monroe_ionphoton_csrbank1_pi0_wrdata2_r;
	end
	if (monroe_ionphoton_csrbank1_pi0_wrdata1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[15:8] <= monroe_ionphoton_csrbank1_pi0_wrdata1_r;
	end
	if (monroe_ionphoton_csrbank1_pi0_wrdata0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi0_wrdata0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_re <= monroe_ionphoton_csrbank1_pi0_wrdata0_re;
	if (monroe_ionphoton_csrbank1_pi1_command0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage_full[5:0] <= monroe_ionphoton_csrbank1_pi1_command0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_re <= monroe_ionphoton_csrbank1_pi1_command0_re;
	if (monroe_ionphoton_csrbank1_pi1_address1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full[14:8] <= monroe_ionphoton_csrbank1_pi1_address1_r;
	end
	if (monroe_ionphoton_csrbank1_pi1_address0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi1_address0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_re <= monroe_ionphoton_csrbank1_pi1_address0_re;
	if (monroe_ionphoton_csrbank1_pi1_baddress0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage_full[2:0] <= monroe_ionphoton_csrbank1_pi1_baddress0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_re <= monroe_ionphoton_csrbank1_pi1_baddress0_re;
	if (monroe_ionphoton_csrbank1_pi1_wrdata3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[31:24] <= monroe_ionphoton_csrbank1_pi1_wrdata3_r;
	end
	if (monroe_ionphoton_csrbank1_pi1_wrdata2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[23:16] <= monroe_ionphoton_csrbank1_pi1_wrdata2_r;
	end
	if (monroe_ionphoton_csrbank1_pi1_wrdata1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[15:8] <= monroe_ionphoton_csrbank1_pi1_wrdata1_r;
	end
	if (monroe_ionphoton_csrbank1_pi1_wrdata0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi1_wrdata0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_re <= monroe_ionphoton_csrbank1_pi1_wrdata0_re;
	if (monroe_ionphoton_csrbank1_pi2_command0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage_full[5:0] <= monroe_ionphoton_csrbank1_pi2_command0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_re <= monroe_ionphoton_csrbank1_pi2_command0_re;
	if (monroe_ionphoton_csrbank1_pi2_address1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full[14:8] <= monroe_ionphoton_csrbank1_pi2_address1_r;
	end
	if (monroe_ionphoton_csrbank1_pi2_address0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi2_address0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_re <= monroe_ionphoton_csrbank1_pi2_address0_re;
	if (monroe_ionphoton_csrbank1_pi2_baddress0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage_full[2:0] <= monroe_ionphoton_csrbank1_pi2_baddress0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_re <= monroe_ionphoton_csrbank1_pi2_baddress0_re;
	if (monroe_ionphoton_csrbank1_pi2_wrdata3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[31:24] <= monroe_ionphoton_csrbank1_pi2_wrdata3_r;
	end
	if (monroe_ionphoton_csrbank1_pi2_wrdata2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[23:16] <= monroe_ionphoton_csrbank1_pi2_wrdata2_r;
	end
	if (monroe_ionphoton_csrbank1_pi2_wrdata1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[15:8] <= monroe_ionphoton_csrbank1_pi2_wrdata1_r;
	end
	if (monroe_ionphoton_csrbank1_pi2_wrdata0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi2_wrdata0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_re <= monroe_ionphoton_csrbank1_pi2_wrdata0_re;
	if (monroe_ionphoton_csrbank1_pi3_command0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage_full[5:0] <= monroe_ionphoton_csrbank1_pi3_command0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_re <= monroe_ionphoton_csrbank1_pi3_command0_re;
	if (monroe_ionphoton_csrbank1_pi3_address1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full[14:8] <= monroe_ionphoton_csrbank1_pi3_address1_r;
	end
	if (monroe_ionphoton_csrbank1_pi3_address0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi3_address0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_re <= monroe_ionphoton_csrbank1_pi3_address0_re;
	if (monroe_ionphoton_csrbank1_pi3_baddress0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage_full[2:0] <= monroe_ionphoton_csrbank1_pi3_baddress0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_re <= monroe_ionphoton_csrbank1_pi3_baddress0_re;
	if (monroe_ionphoton_csrbank1_pi3_wrdata3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[31:24] <= monroe_ionphoton_csrbank1_pi3_wrdata3_r;
	end
	if (monroe_ionphoton_csrbank1_pi3_wrdata2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[23:16] <= monroe_ionphoton_csrbank1_pi3_wrdata2_r;
	end
	if (monroe_ionphoton_csrbank1_pi3_wrdata1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[15:8] <= monroe_ionphoton_csrbank1_pi3_wrdata1_r;
	end
	if (monroe_ionphoton_csrbank1_pi3_wrdata0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full[7:0] <= monroe_ionphoton_csrbank1_pi3_wrdata0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_re <= monroe_ionphoton_csrbank1_pi3_wrdata0_re;
	monroe_ionphoton_interface2_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank2_sel) begin
		case (monroe_ionphoton_interface2_bank_bus_adr[4:0])
			1'd0: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_slot_w;
			end
			1'd1: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_length3_w;
			end
			2'd2: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_length2_w;
			end
			2'd3: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_length1_w;
			end
			3'd4: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_length0_w;
			end
			3'd5: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_errors3_w;
			end
			3'd6: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_errors2_w;
			end
			3'd7: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_errors1_w;
			end
			4'd8: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_errors0_w;
			end
			4'd9: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_writer_status_w;
			end
			4'd10: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_writer_pending_w;
			end
			4'd11: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_writer_ev_enable0_w;
			end
			4'd12: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_reader_start_w;
			end
			4'd13: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_reader_ready_w;
			end
			4'd14: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_reader_slot0_w;
			end
			4'd15: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_reader_length1_w;
			end
			5'd16: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_reader_length0_w;
			end
			5'd17: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_reader_eventmanager_status_w;
			end
			5'd18: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_reader_eventmanager_pending_w;
			end
			5'd19: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_sram_reader_ev_enable0_w;
			end
			5'd20: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_preamble_errors3_w;
			end
			5'd21: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_preamble_errors2_w;
			end
			5'd22: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_preamble_errors1_w;
			end
			5'd23: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_preamble_errors0_w;
			end
			5'd24: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_crc_errors3_w;
			end
			5'd25: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_crc_errors2_w;
			end
			5'd26: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_crc_errors1_w;
			end
			5'd27: begin
				monroe_ionphoton_interface2_bank_bus_dat_r <= monroe_ionphoton_csrbank2_crc_errors0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank2_sram_writer_ev_enable0_re) begin
		monroe_ionphoton_monroe_ionphoton_writer_storage_full <= monroe_ionphoton_csrbank2_sram_writer_ev_enable0_r;
	end
	monroe_ionphoton_monroe_ionphoton_writer_re <= monroe_ionphoton_csrbank2_sram_writer_ev_enable0_re;
	if (monroe_ionphoton_csrbank2_sram_reader_slot0_re) begin
		monroe_ionphoton_monroe_ionphoton_reader_slot_storage_full[1:0] <= monroe_ionphoton_csrbank2_sram_reader_slot0_r;
	end
	monroe_ionphoton_monroe_ionphoton_reader_slot_re <= monroe_ionphoton_csrbank2_sram_reader_slot0_re;
	if (monroe_ionphoton_csrbank2_sram_reader_length1_re) begin
		monroe_ionphoton_monroe_ionphoton_reader_length_storage_full[10:8] <= monroe_ionphoton_csrbank2_sram_reader_length1_r;
	end
	if (monroe_ionphoton_csrbank2_sram_reader_length0_re) begin
		monroe_ionphoton_monroe_ionphoton_reader_length_storage_full[7:0] <= monroe_ionphoton_csrbank2_sram_reader_length0_r;
	end
	monroe_ionphoton_monroe_ionphoton_reader_length_re <= monroe_ionphoton_csrbank2_sram_reader_length0_re;
	if (monroe_ionphoton_csrbank2_sram_reader_ev_enable0_re) begin
		monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage_full <= monroe_ionphoton_csrbank2_sram_reader_ev_enable0_r;
	end
	monroe_ionphoton_monroe_ionphoton_reader_eventmanager_re <= monroe_ionphoton_csrbank2_sram_reader_ev_enable0_re;
	monroe_ionphoton_interface3_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank3_sel) begin
		case (monroe_ionphoton_interface3_bank_bus_adr[1:0])
			1'd0: begin
				monroe_ionphoton_interface3_bank_bus_dat_r <= monroe_ionphoton_csrbank3_in_w;
			end
			1'd1: begin
				monroe_ionphoton_interface3_bank_bus_dat_r <= monroe_ionphoton_csrbank3_out0_w;
			end
			2'd2: begin
				monroe_ionphoton_interface3_bank_bus_dat_r <= monroe_ionphoton_csrbank3_oe0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank3_out0_re) begin
		monroe_ionphoton_i2c_out_storage_full[1:0] <= monroe_ionphoton_csrbank3_out0_r;
	end
	monroe_ionphoton_i2c_out_re <= monroe_ionphoton_csrbank3_out0_re;
	if (monroe_ionphoton_csrbank3_oe0_re) begin
		monroe_ionphoton_i2c_oe_storage_full[1:0] <= monroe_ionphoton_csrbank3_oe0_r;
	end
	monroe_ionphoton_i2c_oe_re <= monroe_ionphoton_csrbank3_oe0_re;
	monroe_ionphoton_interface4_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank4_sel) begin
		case (monroe_ionphoton_interface4_bank_bus_adr[0])
			1'd0: begin
				monroe_ionphoton_interface4_bank_bus_dat_r <= monroe_ionphoton_csrbank4_address0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface4_bank_bus_dat_r <= monroe_ionphoton_csrbank4_data_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank4_address0_re) begin
		monroe_ionphoton_add_identifier_storage_full[7:0] <= monroe_ionphoton_csrbank4_address0_r;
	end
	monroe_ionphoton_add_identifier_re <= monroe_ionphoton_csrbank4_address0_re;
	monroe_ionphoton_interface5_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank5_sel) begin
		case (monroe_ionphoton_interface5_bank_bus_adr[0])
			1'd0: begin
				monroe_ionphoton_interface5_bank_bus_dat_r <= monroe_ionphoton_csrbank5_reset0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank5_reset0_re) begin
		monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage_full <= monroe_ionphoton_csrbank5_reset0_r;
	end
	monroe_ionphoton_monroe_ionphoton_kernel_cpu_re <= monroe_ionphoton_csrbank5_reset0_re;
	monroe_ionphoton_interface6_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank6_sel) begin
		case (monroe_ionphoton_interface6_bank_bus_adr[0])
			1'd0: begin
				monroe_ionphoton_interface6_bank_bus_dat_r <= monroe_ionphoton_csrbank6_out0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank6_out0_re) begin
		monroe_ionphoton_leds_storage_full <= monroe_ionphoton_csrbank6_out0_r;
	end
	monroe_ionphoton_leds_re <= monroe_ionphoton_csrbank6_out0_re;
	monroe_ionphoton_interface7_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank7_sel) begin
		case (monroe_ionphoton_interface7_bank_bus_adr[4:0])
			1'd0: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_enable0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_busy_w;
			end
			2'd2: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_message_encoder_overflow_w;
			end
			2'd3: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_rtio_analyzer_message_encoder_overflow_reset_w;
			end
			3'd4: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_rtio_analyzer_dma_reset_w;
			end
			3'd5: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_base_address4_w;
			end
			3'd6: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_base_address3_w;
			end
			3'd7: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_base_address2_w;
			end
			4'd8: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_base_address1_w;
			end
			4'd9: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_base_address0_w;
			end
			4'd10: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_last_address4_w;
			end
			4'd11: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_last_address3_w;
			end
			4'd12: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_last_address2_w;
			end
			4'd13: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_last_address1_w;
			end
			4'd14: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_last_address0_w;
			end
			4'd15: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count7_w;
			end
			5'd16: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count6_w;
			end
			5'd17: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count5_w;
			end
			5'd18: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count4_w;
			end
			5'd19: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count3_w;
			end
			5'd20: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count2_w;
			end
			5'd21: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count1_w;
			end
			5'd22: begin
				monroe_ionphoton_interface7_bank_bus_dat_r <= monroe_ionphoton_csrbank7_dma_byte_count0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank7_enable0_re) begin
		monroe_ionphoton_rtio_analyzer_enable_storage_full <= monroe_ionphoton_csrbank7_enable0_r;
	end
	monroe_ionphoton_rtio_analyzer_enable_re <= monroe_ionphoton_csrbank7_enable0_re;
	if (monroe_ionphoton_csrbank7_dma_base_address4_re) begin
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[33:32] <= monroe_ionphoton_csrbank7_dma_base_address4_r;
	end
	if (monroe_ionphoton_csrbank7_dma_base_address3_re) begin
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[31:24] <= monroe_ionphoton_csrbank7_dma_base_address3_r;
	end
	if (monroe_ionphoton_csrbank7_dma_base_address2_re) begin
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[23:16] <= monroe_ionphoton_csrbank7_dma_base_address2_r;
	end
	if (monroe_ionphoton_csrbank7_dma_base_address1_re) begin
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[15:8] <= monroe_ionphoton_csrbank7_dma_base_address1_r;
	end
	if (monroe_ionphoton_csrbank7_dma_base_address0_re) begin
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full[7:0] <= monroe_ionphoton_csrbank7_dma_base_address0_r;
	end
	monroe_ionphoton_rtio_analyzer_dma_base_address_re <= monroe_ionphoton_csrbank7_dma_base_address0_re;
	if (monroe_ionphoton_csrbank7_dma_last_address4_re) begin
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[33:32] <= monroe_ionphoton_csrbank7_dma_last_address4_r;
	end
	if (monroe_ionphoton_csrbank7_dma_last_address3_re) begin
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[31:24] <= monroe_ionphoton_csrbank7_dma_last_address3_r;
	end
	if (monroe_ionphoton_csrbank7_dma_last_address2_re) begin
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[23:16] <= monroe_ionphoton_csrbank7_dma_last_address2_r;
	end
	if (monroe_ionphoton_csrbank7_dma_last_address1_re) begin
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[15:8] <= monroe_ionphoton_csrbank7_dma_last_address1_r;
	end
	if (monroe_ionphoton_csrbank7_dma_last_address0_re) begin
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full[7:0] <= monroe_ionphoton_csrbank7_dma_last_address0_r;
	end
	monroe_ionphoton_rtio_analyzer_dma_last_address_re <= monroe_ionphoton_csrbank7_dma_last_address0_re;
	monroe_ionphoton_interface8_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank8_sel) begin
		case (monroe_ionphoton_interface8_bank_bus_adr[3:0])
			1'd0: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_rtio_core_reset_w;
			end
			1'd1: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_rtio_core_reset_phy_w;
			end
			2'd2: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_rtio_core_async_error_w;
			end
			2'd3: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_collision_channel1_w;
			end
			3'd4: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_collision_channel0_w;
			end
			3'd5: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_busy_channel1_w;
			end
			3'd6: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_busy_channel0_w;
			end
			3'd7: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_sequence_error_channel1_w;
			end
			4'd8: begin
				monroe_ionphoton_interface8_bank_bus_dat_r <= monroe_ionphoton_csrbank8_sequence_error_channel0_w;
			end
		endcase
	end
	monroe_ionphoton_interface9_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank9_sel) begin
		case (monroe_ionphoton_interface9_bank_bus_adr[0])
			1'd0: begin
				monroe_ionphoton_interface9_bank_bus_dat_r <= monroe_ionphoton_csrbank9_pll_reset0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface9_bank_bus_dat_r <= monroe_ionphoton_csrbank9_pll_locked_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank9_pll_reset0_re) begin
		monroe_ionphoton_rtio_crg_storage_full <= monroe_ionphoton_csrbank9_pll_reset0_r;
	end
	monroe_ionphoton_rtio_crg_re <= monroe_ionphoton_csrbank9_pll_reset0_re;
	monroe_ionphoton_interface10_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank10_sel) begin
		case (monroe_ionphoton_interface10_bank_bus_adr[2:0])
			1'd0: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_csrbank10_mon_chan_sel0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_csrbank10_mon_probe_sel0_w;
			end
			2'd2: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_mon_value_update_w;
			end
			2'd3: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_csrbank10_mon_value_w;
			end
			3'd4: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_csrbank10_inj_chan_sel0_w;
			end
			3'd5: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_csrbank10_inj_override_sel0_w;
			end
			3'd6: begin
				monroe_ionphoton_interface10_bank_bus_dat_r <= monroe_ionphoton_inj_value_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank10_mon_chan_sel0_re) begin
		monroe_ionphoton_mon_chan_sel_storage_full[5:0] <= monroe_ionphoton_csrbank10_mon_chan_sel0_r;
	end
	monroe_ionphoton_mon_chan_sel_re <= monroe_ionphoton_csrbank10_mon_chan_sel0_re;
	if (monroe_ionphoton_csrbank10_mon_probe_sel0_re) begin
		monroe_ionphoton_mon_probe_sel_storage_full <= monroe_ionphoton_csrbank10_mon_probe_sel0_r;
	end
	monroe_ionphoton_mon_probe_sel_re <= monroe_ionphoton_csrbank10_mon_probe_sel0_re;
	if (monroe_ionphoton_csrbank10_inj_chan_sel0_re) begin
		monroe_ionphoton_inj_chan_sel_storage_full[5:0] <= monroe_ionphoton_csrbank10_inj_chan_sel0_r;
	end
	monroe_ionphoton_inj_chan_sel_re <= monroe_ionphoton_csrbank10_inj_chan_sel0_re;
	if (monroe_ionphoton_csrbank10_inj_override_sel0_re) begin
		monroe_ionphoton_inj_override_sel_storage_full[1:0] <= monroe_ionphoton_csrbank10_inj_override_sel0_r;
	end
	monroe_ionphoton_inj_override_sel_re <= monroe_ionphoton_csrbank10_inj_override_sel0_re;
	monroe_ionphoton_interface11_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank11_sel) begin
		case (monroe_ionphoton_interface11_bank_bus_adr[1:0])
			1'd0: begin
				monroe_ionphoton_interface11_bank_bus_dat_r <= monroe_ionphoton_csrbank11_bitbang0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface11_bank_bus_dat_r <= monroe_ionphoton_csrbank11_miso_w;
			end
			2'd2: begin
				monroe_ionphoton_interface11_bank_bus_dat_r <= monroe_ionphoton_csrbank11_bitbang_en0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank11_bitbang0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage_full[3:0] <= monroe_ionphoton_csrbank11_bitbang0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_re <= monroe_ionphoton_csrbank11_bitbang0_re;
	if (monroe_ionphoton_csrbank11_bitbang_en0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage_full <= monroe_ionphoton_csrbank11_bitbang_en0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_re <= monroe_ionphoton_csrbank11_bitbang_en0_re;
	monroe_ionphoton_interface12_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank12_sel) begin
		case (monroe_ionphoton_interface12_bank_bus_adr[4:0])
			1'd0: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load7_w;
			end
			1'd1: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load6_w;
			end
			2'd2: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load5_w;
			end
			2'd3: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load4_w;
			end
			3'd4: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load3_w;
			end
			3'd5: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load2_w;
			end
			3'd6: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load1_w;
			end
			3'd7: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_load0_w;
			end
			4'd8: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload7_w;
			end
			4'd9: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload6_w;
			end
			4'd10: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload5_w;
			end
			4'd11: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload4_w;
			end
			4'd12: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload3_w;
			end
			4'd13: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload2_w;
			end
			4'd14: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload1_w;
			end
			4'd15: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_reload0_w;
			end
			5'd16: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_en0_w;
			end
			5'd17: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_update_value_w;
			end
			5'd18: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value7_w;
			end
			5'd19: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value6_w;
			end
			5'd20: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value5_w;
			end
			5'd21: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value4_w;
			end
			5'd22: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value3_w;
			end
			5'd23: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value2_w;
			end
			5'd24: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value1_w;
			end
			5'd25: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_value0_w;
			end
			5'd26: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_status_w;
			end
			5'd27: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_pending_w;
			end
			5'd28: begin
				monroe_ionphoton_interface12_bank_bus_dat_r <= monroe_ionphoton_csrbank12_ev_enable0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank12_load7_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[63:56] <= monroe_ionphoton_csrbank12_load7_r;
	end
	if (monroe_ionphoton_csrbank12_load6_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[55:48] <= monroe_ionphoton_csrbank12_load6_r;
	end
	if (monroe_ionphoton_csrbank12_load5_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[47:40] <= monroe_ionphoton_csrbank12_load5_r;
	end
	if (monroe_ionphoton_csrbank12_load4_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[39:32] <= monroe_ionphoton_csrbank12_load4_r;
	end
	if (monroe_ionphoton_csrbank12_load3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[31:24] <= monroe_ionphoton_csrbank12_load3_r;
	end
	if (monroe_ionphoton_csrbank12_load2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[23:16] <= monroe_ionphoton_csrbank12_load2_r;
	end
	if (monroe_ionphoton_csrbank12_load1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[15:8] <= monroe_ionphoton_csrbank12_load1_r;
	end
	if (monroe_ionphoton_csrbank12_load0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full[7:0] <= monroe_ionphoton_csrbank12_load0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_re <= monroe_ionphoton_csrbank12_load0_re;
	if (monroe_ionphoton_csrbank12_reload7_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[63:56] <= monroe_ionphoton_csrbank12_reload7_r;
	end
	if (monroe_ionphoton_csrbank12_reload6_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[55:48] <= monroe_ionphoton_csrbank12_reload6_r;
	end
	if (monroe_ionphoton_csrbank12_reload5_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[47:40] <= monroe_ionphoton_csrbank12_reload5_r;
	end
	if (monroe_ionphoton_csrbank12_reload4_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[39:32] <= monroe_ionphoton_csrbank12_reload4_r;
	end
	if (monroe_ionphoton_csrbank12_reload3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[31:24] <= monroe_ionphoton_csrbank12_reload3_r;
	end
	if (monroe_ionphoton_csrbank12_reload2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[23:16] <= monroe_ionphoton_csrbank12_reload2_r;
	end
	if (monroe_ionphoton_csrbank12_reload1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[15:8] <= monroe_ionphoton_csrbank12_reload1_r;
	end
	if (monroe_ionphoton_csrbank12_reload0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full[7:0] <= monroe_ionphoton_csrbank12_reload0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_re <= monroe_ionphoton_csrbank12_reload0_re;
	if (monroe_ionphoton_csrbank12_en0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage_full <= monroe_ionphoton_csrbank12_en0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_re <= monroe_ionphoton_csrbank12_en0_re;
	if (monroe_ionphoton_csrbank12_ev_enable0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage_full <= monroe_ionphoton_csrbank12_ev_enable0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_re <= monroe_ionphoton_csrbank12_ev_enable0_re;
	monroe_ionphoton_interface13_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank13_sel) begin
		case (monroe_ionphoton_interface13_bank_bus_adr[2:0])
			1'd0: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_enable_null0_w;
			end
			1'd1: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_enable_prog0_w;
			end
			2'd2: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_prog_address3_w;
			end
			2'd3: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_prog_address2_w;
			end
			3'd4: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_prog_address1_w;
			end
			3'd5: begin
				monroe_ionphoton_interface13_bank_bus_dat_r <= monroe_ionphoton_csrbank13_prog_address0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank13_enable_null0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage_full <= monroe_ionphoton_csrbank13_enable_null0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_re <= monroe_ionphoton_csrbank13_enable_null0_re;
	if (monroe_ionphoton_csrbank13_enable_prog0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage_full <= monroe_ionphoton_csrbank13_enable_prog0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_re <= monroe_ionphoton_csrbank13_enable_prog0_re;
	if (monroe_ionphoton_csrbank13_prog_address3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[29:24] <= monroe_ionphoton_csrbank13_prog_address3_r;
	end
	if (monroe_ionphoton_csrbank13_prog_address2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[23:16] <= monroe_ionphoton_csrbank13_prog_address2_r;
	end
	if (monroe_ionphoton_csrbank13_prog_address1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[15:8] <= monroe_ionphoton_csrbank13_prog_address1_r;
	end
	if (monroe_ionphoton_csrbank13_prog_address0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full[7:0] <= monroe_ionphoton_csrbank13_prog_address0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_re <= monroe_ionphoton_csrbank13_prog_address0_re;
	monroe_ionphoton_interface14_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank14_sel) begin
		case (monroe_ionphoton_interface14_bank_bus_adr[2:0])
			1'd0: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rxtx_w;
			end
			1'd1: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_csrbank14_txfull_w;
			end
			2'd2: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_csrbank14_rxempty_w;
			end
			2'd3: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_status_w;
			end
			3'd4: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_pending_w;
			end
			3'd5: begin
				monroe_ionphoton_interface14_bank_bus_dat_r <= monroe_ionphoton_csrbank14_ev_enable0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank14_ev_enable0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage_full[1:0] <= monroe_ionphoton_csrbank14_ev_enable0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_re <= monroe_ionphoton_csrbank14_ev_enable0_re;
	monroe_ionphoton_interface15_bank_bus_dat_r <= 1'd0;
	if (monroe_ionphoton_csrbank15_sel) begin
		case (monroe_ionphoton_interface15_bank_bus_adr[1:0])
			1'd0: begin
				monroe_ionphoton_interface15_bank_bus_dat_r <= monroe_ionphoton_csrbank15_tuning_word3_w;
			end
			1'd1: begin
				monroe_ionphoton_interface15_bank_bus_dat_r <= monroe_ionphoton_csrbank15_tuning_word2_w;
			end
			2'd2: begin
				monroe_ionphoton_interface15_bank_bus_dat_r <= monroe_ionphoton_csrbank15_tuning_word1_w;
			end
			2'd3: begin
				monroe_ionphoton_interface15_bank_bus_dat_r <= monroe_ionphoton_csrbank15_tuning_word0_w;
			end
		endcase
	end
	if (monroe_ionphoton_csrbank15_tuning_word3_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[31:24] <= monroe_ionphoton_csrbank15_tuning_word3_r;
	end
	if (monroe_ionphoton_csrbank15_tuning_word2_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[23:16] <= monroe_ionphoton_csrbank15_tuning_word2_r;
	end
	if (monroe_ionphoton_csrbank15_tuning_word1_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[15:8] <= monroe_ionphoton_csrbank15_tuning_word1_r;
	end
	if (monroe_ionphoton_csrbank15_tuning_word0_re) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full[7:0] <= monroe_ionphoton_csrbank15_tuning_word0_r;
	end
	monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_re <= monroe_ionphoton_csrbank15_tuning_word0_re;
	if (sys_rst) begin
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_null_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_enable_prog_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_storage_full <= 30'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_prog_address_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tmpu_error <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_bus_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_adr <= 14'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_we <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interface_dat_w <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_bus_wishbone_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_counter <= 2'd0;
		serial_tx <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_storage_full <= 32'd4367715;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_sink_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_txen <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_tx <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_reg <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_bitcount <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_tx_busy <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_stb <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_source_payload_data <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_uart_clk_rxen <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_phase_accumulator_rx <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_r <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_reg <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_bitcount <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_phy_rx_busy <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_pending <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_old_trigger <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_pending <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_old_trigger <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_storage_full <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_level <= 5'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_produce <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_consume <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_level <= 5'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_produce <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_consume <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_storage_full <= 64'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_load_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_storage_full <= 64'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_reload_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_en_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value_status <= 64'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_pending <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_zero_old_trigger <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_eventmanager_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_timer0_value <= 64'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage_full <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dqs <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en2 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en3 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_n_rddata_en4 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_last_wrdata_en <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_storage_full <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_storage_full <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_command_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_storage_full <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_address_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_storage_full <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_baddress_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_storage_full <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_wrdata_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector0_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_storage_full <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_command_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_storage_full <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_address_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_storage_full <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_baddress_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_storage_full <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_wrdata_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector1_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_storage_full <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_command_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_storage_full <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_address_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_storage_full <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_baddress_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_storage_full <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_wrdata_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector2_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_storage_full <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_command_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_storage_full <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_address_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_storage_full <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_baddress_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_storage_full <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_wrdata_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_phaseinjector3_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank0_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank1_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank2_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank3_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank4_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank5_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank6_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_idle <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_bank7_row1 <= 15'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_write2precharge_timer_count <= 3'd4;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sdram_controller_refresh_timer_count <= 10'd886;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_adr_offset_r <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bus_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_storage_full <= 4'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_bitbang_en_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_cs_n <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_clk <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dq_oe <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_sr <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_dqi <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_counter <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_tx_mmcm_reset <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_rx_mmcm_reset <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_tx_init_qpll_reset0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_tx_init_tx_reset0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_tx_init_timer <= 6'd0;
		monroe_ionphoton_monroe_ionphoton_tx_init_tick <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_rx_init_rx_reset0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_rx_init_drpvalue <= 16'd0;
		monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done_r <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_cdr_lock_counter <= 13'd0;
		monroe_ionphoton_monroe_ionphoton_cdr_locked <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_preamble_errors_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_crc_errors_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter0_q_binary <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter1_q_binary <= 7'd0;
		monroe_ionphoton_monroe_ionphoton_writer_errors_status <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_writer_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_writer_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_writer_counter <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_writer_slot <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_writer_fifo_level <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_writer_fifo_produce <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_writer_fifo_consume <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_reader_slot_storage_full <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_reader_slot_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_reader_length_storage_full <= 11'd0;
		monroe_ionphoton_monroe_ionphoton_reader_length_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_reader_done_pending <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_reader_eventmanager_storage_full <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_reader_eventmanager_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_reader_fifo_level <= 3'd0;
		monroe_ionphoton_monroe_ionphoton_reader_fifo_produce <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_reader_fifo_consume <= 2'd0;
		monroe_ionphoton_monroe_ionphoton_reader_counter <= 11'd0;
		monroe_ionphoton_monroe_ionphoton_reader_last_d <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram0_bus_ack0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram1_bus_ack0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram2_bus_ack0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram3_bus_ack0 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram0_bus_ack1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram1_bus_ack1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram2_bus_ack1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_sram3_bus_ack1 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_slave_sel_r <= 8'd0;
		monroe_ionphoton_monroe_ionphoton_kernel_cpu_storage_full <= 1'd1;
		monroe_ionphoton_monroe_ionphoton_kernel_cpu_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox_i1_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox_i1_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox_i2_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox_i2_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox0 <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox1 <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_mailbox2 <= 32'd0;
		monroe_ionphoton_add_identifier_storage_full <= 8'd0;
		monroe_ionphoton_add_identifier_re <= 1'd0;
		monroe_ionphoton_leds_storage_full <= 1'd0;
		monroe_ionphoton_leds_re <= 1'd0;
		monroe_ionphoton_i2c_out_storage_full <= 2'd0;
		monroe_ionphoton_i2c_out_re <= 1'd0;
		monroe_ionphoton_i2c_oe_storage_full <= 2'd0;
		monroe_ionphoton_i2c_oe_re <= 1'd0;
		monroe_ionphoton_rtio_crg_storage_full <= 1'd1;
		monroe_ionphoton_rtio_crg_re <= 1'd0;
		monroe_ionphoton_rtio_core_collision_channel_status <= 16'd0;
		monroe_ionphoton_rtio_core_busy_channel_status <= 16'd0;
		monroe_ionphoton_rtio_core_sequence_error_channel_status <= 16'd0;
		monroe_ionphoton_rtio_core_cmd_reset <= 1'd1;
		monroe_ionphoton_rtio_core_cmd_reset_phy <= 1'd1;
		monroe_ionphoton_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= 61'd0;
		monroe_ionphoton_rtio_core_o_collision <= 1'd0;
		monroe_ionphoton_rtio_core_o_busy <= 1'd0;
		monroe_ionphoton_rtio_core_o_sequence_error <= 1'd0;
		monroe_ionphoton_rtio_target_storage_full <= 32'd0;
		monroe_ionphoton_rtio_target_re <= 1'd0;
		monroe_ionphoton_rtio_o_data_storage_full <= 512'd0;
		monroe_ionphoton_rtio_o_data_re <= 1'd0;
		monroe_ionphoton_rtio_i_timeout_storage_full <= 64'd0;
		monroe_ionphoton_rtio_i_timeout_re <= 1'd0;
		monroe_ionphoton_rtio_counter_status <= 64'd0;
		monroe_ionphoton_rtio_now_hi_backing <= 32'd0;
		monroe_ionphoton_dma_dma_storage_full <= 34'd0;
		monroe_ionphoton_dma_dma_re <= 1'd0;
		monroe_ionphoton_dma_time_offset_storage_full <= 64'd0;
		monroe_ionphoton_dma_time_offset_re <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank0_bus_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank0_bus_ack <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank1_bus_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank1_bus_ack <= 1'd0;
		monroe_ionphoton_cri_con_storage_full <= 2'd0;
		monroe_ionphoton_cri_con_re <= 1'd0;
		monroe_ionphoton_cri_con_selected <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank2_bus_dat_r <= 32'd0;
		monroe_ionphoton_monroe_ionphoton_csrbank2_bus_ack <= 1'd0;
		monroe_ionphoton_mon_chan_sel_storage_full <= 6'd0;
		monroe_ionphoton_mon_chan_sel_re <= 1'd0;
		monroe_ionphoton_mon_probe_sel_storage_full <= 1'd0;
		monroe_ionphoton_mon_probe_sel_re <= 1'd0;
		monroe_ionphoton_mon_status <= 1'd0;
		monroe_ionphoton_inj_chan_sel_storage_full <= 6'd0;
		monroe_ionphoton_inj_chan_sel_re <= 1'd0;
		monroe_ionphoton_inj_override_sel_storage_full <= 2'd0;
		monroe_ionphoton_inj_override_sel_re <= 1'd0;
		monroe_ionphoton_inj_o_sys0 <= 1'd0;
		monroe_ionphoton_inj_o_sys1 <= 1'd0;
		monroe_ionphoton_inj_o_sys2 <= 1'd0;
		monroe_ionphoton_inj_o_sys3 <= 1'd0;
		monroe_ionphoton_inj_o_sys4 <= 1'd0;
		monroe_ionphoton_inj_o_sys5 <= 1'd0;
		monroe_ionphoton_inj_o_sys6 <= 1'd0;
		monroe_ionphoton_inj_o_sys7 <= 1'd0;
		monroe_ionphoton_inj_o_sys8 <= 1'd0;
		monroe_ionphoton_inj_o_sys9 <= 1'd0;
		monroe_ionphoton_inj_o_sys10 <= 1'd0;
		monroe_ionphoton_inj_o_sys11 <= 1'd0;
		monroe_ionphoton_inj_o_sys12 <= 1'd0;
		monroe_ionphoton_inj_o_sys13 <= 1'd0;
		monroe_ionphoton_inj_o_sys14 <= 1'd0;
		monroe_ionphoton_inj_o_sys15 <= 1'd0;
		monroe_ionphoton_inj_o_sys16 <= 1'd0;
		monroe_ionphoton_inj_o_sys17 <= 1'd0;
		monroe_ionphoton_inj_o_sys18 <= 1'd0;
		monroe_ionphoton_inj_o_sys19 <= 1'd0;
		monroe_ionphoton_inj_o_sys20 <= 1'd0;
		monroe_ionphoton_inj_o_sys21 <= 1'd0;
		monroe_ionphoton_inj_o_sys22 <= 1'd0;
		monroe_ionphoton_inj_o_sys23 <= 1'd0;
		monroe_ionphoton_inj_o_sys24 <= 1'd0;
		monroe_ionphoton_inj_o_sys25 <= 1'd0;
		monroe_ionphoton_inj_o_sys26 <= 1'd0;
		monroe_ionphoton_inj_o_sys27 <= 1'd0;
		monroe_ionphoton_inj_o_sys28 <= 1'd0;
		monroe_ionphoton_inj_o_sys29 <= 1'd0;
		monroe_ionphoton_inj_o_sys30 <= 1'd0;
		monroe_ionphoton_inj_o_sys31 <= 1'd0;
		monroe_ionphoton_inj_o_sys32 <= 1'd0;
		monroe_ionphoton_inj_o_sys33 <= 1'd0;
		monroe_ionphoton_inj_o_sys34 <= 1'd0;
		monroe_ionphoton_inj_o_sys35 <= 1'd0;
		monroe_ionphoton_inj_o_sys36 <= 1'd0;
		monroe_ionphoton_inj_o_sys37 <= 1'd0;
		monroe_ionphoton_inj_o_sys38 <= 1'd0;
		monroe_ionphoton_inj_o_sys39 <= 1'd0;
		monroe_ionphoton_inj_o_sys40 <= 1'd0;
		monroe_ionphoton_inj_o_sys41 <= 1'd0;
		monroe_ionphoton_inj_o_sys42 <= 1'd0;
		monroe_ionphoton_inj_o_sys43 <= 1'd0;
		monroe_ionphoton_inj_o_sys44 <= 1'd0;
		monroe_ionphoton_inj_o_sys45 <= 1'd0;
		monroe_ionphoton_inj_o_sys46 <= 1'd0;
		monroe_ionphoton_inj_o_sys47 <= 1'd0;
		monroe_ionphoton_inj_o_sys48 <= 1'd0;
		monroe_ionphoton_inj_o_sys49 <= 1'd0;
		monroe_ionphoton_inj_o_sys50 <= 1'd0;
		monroe_ionphoton_inj_o_sys51 <= 1'd0;
		monroe_ionphoton_inj_o_sys52 <= 1'd0;
		monroe_ionphoton_inj_o_sys53 <= 1'd0;
		monroe_ionphoton_inj_o_sys54 <= 1'd0;
		monroe_ionphoton_inj_o_sys55 <= 1'd0;
		monroe_ionphoton_inj_o_sys56 <= 1'd0;
		monroe_ionphoton_inj_o_sys57 <= 1'd0;
		monroe_ionphoton_inj_o_sys58 <= 1'd0;
		monroe_ionphoton_inj_o_sys59 <= 1'd0;
		monroe_ionphoton_inj_o_sys60 <= 1'd0;
		monroe_ionphoton_inj_o_sys61 <= 1'd0;
		monroe_ionphoton_inj_o_sys62 <= 1'd0;
		monroe_ionphoton_inj_o_sys63 <= 1'd0;
		monroe_ionphoton_inj_o_sys64 <= 1'd0;
		monroe_ionphoton_inj_o_sys65 <= 1'd0;
		monroe_ionphoton_inj_o_sys66 <= 1'd0;
		monroe_ionphoton_inj_o_sys67 <= 1'd0;
		monroe_ionphoton_inj_o_sys68 <= 1'd0;
		monroe_ionphoton_inj_o_sys69 <= 1'd0;
		monroe_ionphoton_monroe_ionphoton_interface1_bus_adr <= 30'd0;
		monroe_ionphoton_rtio_analyzer_enable_storage_full <= 1'd0;
		monroe_ionphoton_rtio_analyzer_enable_re <= 1'd0;
		monroe_ionphoton_rtio_analyzer_busy_status <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_source_stb <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_source_payload_data <= 256'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_status <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_read_wait_event_r <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_just_written <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_enable_r <= 1'd0;
		monroe_ionphoton_rtio_analyzer_message_encoder_stopping <= 1'd0;
		monroe_ionphoton_rtio_analyzer_fifo_readable <= 1'd0;
		monroe_ionphoton_rtio_analyzer_fifo_level0 <= 8'd0;
		monroe_ionphoton_rtio_analyzer_fifo_produce <= 7'd0;
		monroe_ionphoton_rtio_analyzer_fifo_consume <= 7'd0;
		monroe_ionphoton_rtio_analyzer_converter_mux <= 1'd0;
		monroe_ionphoton_rtio_analyzer_dma_base_address_storage_full <= 34'd0;
		monroe_ionphoton_rtio_analyzer_dma_base_address_re <= 1'd0;
		monroe_ionphoton_rtio_analyzer_dma_last_address_storage_full <= 34'd0;
		monroe_ionphoton_rtio_analyzer_dma_last_address_re <= 1'd0;
		monroe_ionphoton_rtio_analyzer_dma_message_count <= 59'd0;
		monroe_ionphoton_rtio_analyzer_enable_r <= 1'd0;
		minicon_state <= 6'd0;
		fullmemorywe_state <= 3'd0;
		a7_1000basex_gtptxinit_state <= 2'd0;
		a7_1000basex_gtprxinit_state <= 4'd0;
		liteethmacsramwriter_state <= 2'd0;
		liteethmacsramreader_state <= 2'd0;
		grant <= 1'd0;
		slave_sel_r <= 5'd0;
		sdram_cpulevel_arbiter_grant <= 1'd0;
		sdram_native_arbiter_grant <= 2'd0;
		monroe_ionphoton_grant <= 1'd0;
		monroe_ionphoton_slave_sel_r <= 6'd0;
		monroe_ionphoton_interface0_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface1_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface2_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface3_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface4_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface5_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface6_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface7_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface8_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface9_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface10_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface11_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface12_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface13_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface14_bank_bus_dat_r <= 8'd0;
		monroe_ionphoton_interface15_bank_bus_dat_r <= 8'd0;
	end
	xilinxmultiregimpl0_regs0 <= serial_rx;
	xilinxmultiregimpl0_regs1 <= xilinxmultiregimpl0_regs0;
	xilinxmultiregimpl4_regs0 <= monroe_ionphoton_monroe_ionphoton_tx_init_qpll_lock0;
	xilinxmultiregimpl4_regs1 <= xilinxmultiregimpl4_regs0;
	xilinxmultiregimpl5_regs0 <= monroe_ionphoton_monroe_ionphoton_rx_init_rx_pma_reset_done0;
	xilinxmultiregimpl5_regs1 <= xilinxmultiregimpl5_regs0;
	xilinxmultiregimpl6_regs0 <= monroe_ionphoton_monroe_ionphoton_toggle_i;
	xilinxmultiregimpl6_regs1 <= xilinxmultiregimpl6_regs0;
	xilinxmultiregimpl7_regs0 <= monroe_ionphoton_monroe_ionphoton_ps_preamble_error_toggle_i;
	xilinxmultiregimpl7_regs1 <= xilinxmultiregimpl7_regs0;
	xilinxmultiregimpl8_regs0 <= monroe_ionphoton_monroe_ionphoton_ps_crc_error_toggle_i;
	xilinxmultiregimpl8_regs1 <= xilinxmultiregimpl8_regs0;
	xilinxmultiregimpl10_regs0 <= monroe_ionphoton_monroe_ionphoton_tx_cdc_graycounter1_q;
	xilinxmultiregimpl10_regs1 <= xilinxmultiregimpl10_regs0;
	xilinxmultiregimpl11_regs0 <= monroe_ionphoton_monroe_ionphoton_rx_cdc_graycounter0_q;
	xilinxmultiregimpl11_regs1 <= xilinxmultiregimpl11_regs0;
	xilinxmultiregimpl13_regs0 <= monroe_ionphoton_i2c_tstriple0_i;
	xilinxmultiregimpl13_regs1 <= xilinxmultiregimpl13_regs0;
	xilinxmultiregimpl14_regs0 <= monroe_ionphoton_i2c_tstriple1_i;
	xilinxmultiregimpl14_regs1 <= xilinxmultiregimpl14_regs0;
	xilinxmultiregimpl15_regs0 <= monroe_ionphoton_rtio_crg_pll_locked;
	xilinxmultiregimpl15_regs1 <= xilinxmultiregimpl15_regs0;
	xilinxmultiregimpl16_regs0 <= monroe_ionphoton_rtio_tsc_value_gray_rtio;
	xilinxmultiregimpl16_regs1 <= xilinxmultiregimpl16_regs0;
	xilinxmultiregimpl67_regs0 <= monroe_ionphoton_mon_bussynchronizer0_i;
	xilinxmultiregimpl67_regs1 <= xilinxmultiregimpl67_regs0;
	xilinxmultiregimpl68_regs0 <= monroe_ionphoton_mon_bussynchronizer1_i;
	xilinxmultiregimpl68_regs1 <= xilinxmultiregimpl68_regs0;
	xilinxmultiregimpl69_regs0 <= monroe_ionphoton_mon_bussynchronizer2_i;
	xilinxmultiregimpl69_regs1 <= xilinxmultiregimpl69_regs0;
	xilinxmultiregimpl70_regs0 <= monroe_ionphoton_mon_bussynchronizer3_i;
	xilinxmultiregimpl70_regs1 <= xilinxmultiregimpl70_regs0;
	xilinxmultiregimpl71_regs0 <= monroe_ionphoton_mon_bussynchronizer4_i;
	xilinxmultiregimpl71_regs1 <= xilinxmultiregimpl71_regs0;
	xilinxmultiregimpl72_regs0 <= monroe_ionphoton_mon_bussynchronizer5_i;
	xilinxmultiregimpl72_regs1 <= xilinxmultiregimpl72_regs0;
	xilinxmultiregimpl73_regs0 <= monroe_ionphoton_mon_bussynchronizer6_i;
	xilinxmultiregimpl73_regs1 <= xilinxmultiregimpl73_regs0;
	xilinxmultiregimpl74_regs0 <= monroe_ionphoton_mon_bussynchronizer7_i;
	xilinxmultiregimpl74_regs1 <= xilinxmultiregimpl74_regs0;
	xilinxmultiregimpl75_regs0 <= monroe_ionphoton_mon_bussynchronizer8_i;
	xilinxmultiregimpl75_regs1 <= xilinxmultiregimpl75_regs0;
	xilinxmultiregimpl76_regs0 <= monroe_ionphoton_mon_bussynchronizer9_i;
	xilinxmultiregimpl76_regs1 <= xilinxmultiregimpl76_regs0;
	xilinxmultiregimpl77_regs0 <= monroe_ionphoton_mon_bussynchronizer10_i;
	xilinxmultiregimpl77_regs1 <= xilinxmultiregimpl77_regs0;
	xilinxmultiregimpl78_regs0 <= monroe_ionphoton_mon_bussynchronizer11_i;
	xilinxmultiregimpl78_regs1 <= xilinxmultiregimpl78_regs0;
	xilinxmultiregimpl79_regs0 <= monroe_ionphoton_mon_bussynchronizer12_i;
	xilinxmultiregimpl79_regs1 <= xilinxmultiregimpl79_regs0;
	xilinxmultiregimpl80_regs0 <= monroe_ionphoton_mon_bussynchronizer13_i;
	xilinxmultiregimpl80_regs1 <= xilinxmultiregimpl80_regs0;
	xilinxmultiregimpl81_regs0 <= monroe_ionphoton_mon_bussynchronizer14_i;
	xilinxmultiregimpl81_regs1 <= xilinxmultiregimpl81_regs0;
	xilinxmultiregimpl82_regs0 <= monroe_ionphoton_mon_bussynchronizer15_i;
	xilinxmultiregimpl82_regs1 <= xilinxmultiregimpl82_regs0;
	xilinxmultiregimpl83_regs0 <= monroe_ionphoton_mon_bussynchronizer16_i;
	xilinxmultiregimpl83_regs1 <= xilinxmultiregimpl83_regs0;
	xilinxmultiregimpl84_regs0 <= monroe_ionphoton_mon_bussynchronizer17_i;
	xilinxmultiregimpl84_regs1 <= xilinxmultiregimpl84_regs0;
	xilinxmultiregimpl85_regs0 <= monroe_ionphoton_mon_bussynchronizer18_i;
	xilinxmultiregimpl85_regs1 <= xilinxmultiregimpl85_regs0;
	xilinxmultiregimpl86_regs0 <= monroe_ionphoton_mon_bussynchronizer19_i;
	xilinxmultiregimpl86_regs1 <= xilinxmultiregimpl86_regs0;
	xilinxmultiregimpl87_regs0 <= monroe_ionphoton_mon_bussynchronizer20_i;
	xilinxmultiregimpl87_regs1 <= xilinxmultiregimpl87_regs0;
	xilinxmultiregimpl88_regs0 <= monroe_ionphoton_mon_bussynchronizer21_i;
	xilinxmultiregimpl88_regs1 <= xilinxmultiregimpl88_regs0;
	xilinxmultiregimpl89_regs0 <= monroe_ionphoton_mon_bussynchronizer22_i;
	xilinxmultiregimpl89_regs1 <= xilinxmultiregimpl89_regs0;
	xilinxmultiregimpl90_regs0 <= monroe_ionphoton_mon_bussynchronizer23_i;
	xilinxmultiregimpl90_regs1 <= xilinxmultiregimpl90_regs0;
	xilinxmultiregimpl91_regs0 <= monroe_ionphoton_mon_bussynchronizer24_i;
	xilinxmultiregimpl91_regs1 <= xilinxmultiregimpl91_regs0;
	xilinxmultiregimpl92_regs0 <= monroe_ionphoton_mon_bussynchronizer25_i;
	xilinxmultiregimpl92_regs1 <= xilinxmultiregimpl92_regs0;
	xilinxmultiregimpl93_regs0 <= monroe_ionphoton_mon_bussynchronizer26_i;
	xilinxmultiregimpl93_regs1 <= xilinxmultiregimpl93_regs0;
	xilinxmultiregimpl94_regs0 <= monroe_ionphoton_mon_bussynchronizer27_i;
	xilinxmultiregimpl94_regs1 <= xilinxmultiregimpl94_regs0;
	xilinxmultiregimpl95_regs0 <= monroe_ionphoton_mon_bussynchronizer28_i;
	xilinxmultiregimpl95_regs1 <= xilinxmultiregimpl95_regs0;
	xilinxmultiregimpl96_regs0 <= monroe_ionphoton_mon_bussynchronizer29_i;
	xilinxmultiregimpl96_regs1 <= xilinxmultiregimpl96_regs0;
	xilinxmultiregimpl97_regs0 <= monroe_ionphoton_mon_bussynchronizer30_i;
	xilinxmultiregimpl97_regs1 <= xilinxmultiregimpl97_regs0;
	xilinxmultiregimpl98_regs0 <= monroe_ionphoton_mon_bussynchronizer31_i;
	xilinxmultiregimpl98_regs1 <= xilinxmultiregimpl98_regs0;
	xilinxmultiregimpl99_regs0 <= monroe_ionphoton_mon_bussynchronizer32_i;
	xilinxmultiregimpl99_regs1 <= xilinxmultiregimpl99_regs0;
	xilinxmultiregimpl100_regs0 <= monroe_ionphoton_mon_bussynchronizer33_i;
	xilinxmultiregimpl100_regs1 <= xilinxmultiregimpl100_regs0;
	xilinxmultiregimpl101_regs0 <= monroe_ionphoton_mon_bussynchronizer34_i;
	xilinxmultiregimpl101_regs1 <= xilinxmultiregimpl101_regs0;
	xilinxmultiregimpl102_regs0 <= monroe_ionphoton_mon_bussynchronizer35_i;
	xilinxmultiregimpl102_regs1 <= xilinxmultiregimpl102_regs0;
	xilinxmultiregimpl103_regs0 <= monroe_ionphoton_mon_bussynchronizer36_i;
	xilinxmultiregimpl103_regs1 <= xilinxmultiregimpl103_regs0;
end

always @(posedge sys_kernel_clk) begin
	monroe_ionphoton_dma_dma_enable_r <= monroe_ionphoton_dma_flow_enable;
	if ((monroe_ionphoton_dma_flow_enable & (~monroe_ionphoton_dma_dma_enable_r))) begin
		monroe_ionphoton_dma_dma_sink_payload_address <= monroe_ionphoton_dma_dma_storage;
		monroe_ionphoton_dma_dma_sink_eop <= 1'd0;
		monroe_ionphoton_dma_dma_sink_stb <= 1'd1;
	end
	if ((monroe_ionphoton_dma_dma_sink_stb & monroe_ionphoton_dma_dma_sink_ack)) begin
		if (monroe_ionphoton_dma_dma_sink_eop) begin
			monroe_ionphoton_dma_dma_sink_stb <= 1'd0;
		end else begin
			monroe_ionphoton_dma_dma_sink_payload_address <= (monroe_ionphoton_dma_dma_sink_payload_address + 1'd1);
			if ((~monroe_ionphoton_dma_flow_enable)) begin
				monroe_ionphoton_dma_dma_sink_eop <= 1'd1;
			end
		end
	end
	if (monroe_ionphoton_dma_dma_source_ack) begin
		monroe_ionphoton_dma_dma_data_reg_loaded <= 1'd0;
	end
	if (monroe_ionphoton_monroe_ionphoton_interface0_bus_ack) begin
		monroe_ionphoton_dma_dma_data_reg_loaded <= 1'd1;
		monroe_ionphoton_dma_dma_source_payload_data <= monroe_ionphoton_monroe_ionphoton_interface0_bus_dat_r;
		monroe_ionphoton_dma_dma_source_eop <= monroe_ionphoton_dma_dma_sink_eop;
	end
	monroe_ionphoton_dma_rawslicer_level <= monroe_ionphoton_dma_rawslicer_next_level;
	if (monroe_ionphoton_dma_rawslicer_load_buf) begin
		case (monroe_ionphoton_dma_rawslicer_level)
			1'd0: begin
				monroe_ionphoton_dma_rawslicer_buf[127:0] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			1'd1: begin
				monroe_ionphoton_dma_rawslicer_buf[135:8] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd2: begin
				monroe_ionphoton_dma_rawslicer_buf[143:16] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			2'd3: begin
				monroe_ionphoton_dma_rawslicer_buf[151:24] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd4: begin
				monroe_ionphoton_dma_rawslicer_buf[159:32] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd5: begin
				monroe_ionphoton_dma_rawslicer_buf[167:40] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd6: begin
				monroe_ionphoton_dma_rawslicer_buf[175:48] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			3'd7: begin
				monroe_ionphoton_dma_rawslicer_buf[183:56] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd8: begin
				monroe_ionphoton_dma_rawslicer_buf[191:64] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd9: begin
				monroe_ionphoton_dma_rawslicer_buf[199:72] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd10: begin
				monroe_ionphoton_dma_rawslicer_buf[207:80] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd11: begin
				monroe_ionphoton_dma_rawslicer_buf[215:88] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd12: begin
				monroe_ionphoton_dma_rawslicer_buf[223:96] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd13: begin
				monroe_ionphoton_dma_rawslicer_buf[231:104] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd14: begin
				monroe_ionphoton_dma_rawslicer_buf[239:112] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			4'd15: begin
				monroe_ionphoton_dma_rawslicer_buf[247:120] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd16: begin
				monroe_ionphoton_dma_rawslicer_buf[255:128] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd17: begin
				monroe_ionphoton_dma_rawslicer_buf[263:136] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd18: begin
				monroe_ionphoton_dma_rawslicer_buf[271:144] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd19: begin
				monroe_ionphoton_dma_rawslicer_buf[279:152] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd20: begin
				monroe_ionphoton_dma_rawslicer_buf[287:160] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd21: begin
				monroe_ionphoton_dma_rawslicer_buf[295:168] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd22: begin
				monroe_ionphoton_dma_rawslicer_buf[303:176] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd23: begin
				monroe_ionphoton_dma_rawslicer_buf[311:184] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd24: begin
				monroe_ionphoton_dma_rawslicer_buf[319:192] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd25: begin
				monroe_ionphoton_dma_rawslicer_buf[327:200] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd26: begin
				monroe_ionphoton_dma_rawslicer_buf[335:208] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd27: begin
				monroe_ionphoton_dma_rawslicer_buf[343:216] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd28: begin
				monroe_ionphoton_dma_rawslicer_buf[351:224] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd29: begin
				monroe_ionphoton_dma_rawslicer_buf[359:232] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd30: begin
				monroe_ionphoton_dma_rawslicer_buf[367:240] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			5'd31: begin
				monroe_ionphoton_dma_rawslicer_buf[375:248] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd32: begin
				monroe_ionphoton_dma_rawslicer_buf[383:256] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd33: begin
				monroe_ionphoton_dma_rawslicer_buf[391:264] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd34: begin
				monroe_ionphoton_dma_rawslicer_buf[399:272] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd35: begin
				monroe_ionphoton_dma_rawslicer_buf[407:280] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd36: begin
				monroe_ionphoton_dma_rawslicer_buf[415:288] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd37: begin
				monroe_ionphoton_dma_rawslicer_buf[423:296] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd38: begin
				monroe_ionphoton_dma_rawslicer_buf[431:304] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd39: begin
				monroe_ionphoton_dma_rawslicer_buf[439:312] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd40: begin
				monroe_ionphoton_dma_rawslicer_buf[447:320] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd41: begin
				monroe_ionphoton_dma_rawslicer_buf[455:328] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd42: begin
				monroe_ionphoton_dma_rawslicer_buf[463:336] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd43: begin
				monroe_ionphoton_dma_rawslicer_buf[471:344] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd44: begin
				monroe_ionphoton_dma_rawslicer_buf[479:352] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd45: begin
				monroe_ionphoton_dma_rawslicer_buf[487:360] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd46: begin
				monroe_ionphoton_dma_rawslicer_buf[495:368] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd47: begin
				monroe_ionphoton_dma_rawslicer_buf[503:376] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd48: begin
				monroe_ionphoton_dma_rawslicer_buf[511:384] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd49: begin
				monroe_ionphoton_dma_rawslicer_buf[519:392] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd50: begin
				monroe_ionphoton_dma_rawslicer_buf[527:400] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd51: begin
				monroe_ionphoton_dma_rawslicer_buf[535:408] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd52: begin
				monroe_ionphoton_dma_rawslicer_buf[543:416] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd53: begin
				monroe_ionphoton_dma_rawslicer_buf[551:424] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd54: begin
				monroe_ionphoton_dma_rawslicer_buf[559:432] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd55: begin
				monroe_ionphoton_dma_rawslicer_buf[567:440] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd56: begin
				monroe_ionphoton_dma_rawslicer_buf[575:448] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd57: begin
				monroe_ionphoton_dma_rawslicer_buf[583:456] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd58: begin
				monroe_ionphoton_dma_rawslicer_buf[591:464] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd59: begin
				monroe_ionphoton_dma_rawslicer_buf[599:472] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd60: begin
				monroe_ionphoton_dma_rawslicer_buf[607:480] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd61: begin
				monroe_ionphoton_dma_rawslicer_buf[615:488] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd62: begin
				monroe_ionphoton_dma_rawslicer_buf[623:496] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			6'd63: begin
				monroe_ionphoton_dma_rawslicer_buf[631:504] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd64: begin
				monroe_ionphoton_dma_rawslicer_buf[639:512] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd65: begin
				monroe_ionphoton_dma_rawslicer_buf[647:520] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd66: begin
				monroe_ionphoton_dma_rawslicer_buf[655:528] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd67: begin
				monroe_ionphoton_dma_rawslicer_buf[663:536] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd68: begin
				monroe_ionphoton_dma_rawslicer_buf[671:544] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd69: begin
				monroe_ionphoton_dma_rawslicer_buf[679:552] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd70: begin
				monroe_ionphoton_dma_rawslicer_buf[687:560] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd71: begin
				monroe_ionphoton_dma_rawslicer_buf[695:568] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd72: begin
				monroe_ionphoton_dma_rawslicer_buf[703:576] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd73: begin
				monroe_ionphoton_dma_rawslicer_buf[711:584] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd74: begin
				monroe_ionphoton_dma_rawslicer_buf[719:592] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd75: begin
				monroe_ionphoton_dma_rawslicer_buf[727:600] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
			7'd76: begin
				monroe_ionphoton_dma_rawslicer_buf[735:608] <= {monroe_ionphoton_dma_rawslicer_sink_payload_data[7:0], monroe_ionphoton_dma_rawslicer_sink_payload_data[15:8], monroe_ionphoton_dma_rawslicer_sink_payload_data[23:16], monroe_ionphoton_dma_rawslicer_sink_payload_data[31:24], monroe_ionphoton_dma_rawslicer_sink_payload_data[39:32], monroe_ionphoton_dma_rawslicer_sink_payload_data[47:40], monroe_ionphoton_dma_rawslicer_sink_payload_data[55:48], monroe_ionphoton_dma_rawslicer_sink_payload_data[63:56], monroe_ionphoton_dma_rawslicer_sink_payload_data[71:64], monroe_ionphoton_dma_rawslicer_sink_payload_data[79:72], monroe_ionphoton_dma_rawslicer_sink_payload_data[87:80], monroe_ionphoton_dma_rawslicer_sink_payload_data[95:88], monroe_ionphoton_dma_rawslicer_sink_payload_data[103:96], monroe_ionphoton_dma_rawslicer_sink_payload_data[111:104], monroe_ionphoton_dma_rawslicer_sink_payload_data[119:112], monroe_ionphoton_dma_rawslicer_sink_payload_data[127:120]};
			end
		endcase
	end
	if (monroe_ionphoton_dma_rawslicer_shift_buf) begin
		case (monroe_ionphoton_dma_rawslicer_source_consume)
			1'd0: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:0];
			end
			1'd1: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:8];
			end
			2'd2: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:16];
			end
			2'd3: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:24];
			end
			3'd4: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:32];
			end
			3'd5: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:40];
			end
			3'd6: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:48];
			end
			3'd7: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:56];
			end
			4'd8: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:64];
			end
			4'd9: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:72];
			end
			4'd10: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:80];
			end
			4'd11: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:88];
			end
			4'd12: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:96];
			end
			4'd13: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:104];
			end
			4'd14: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:112];
			end
			4'd15: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:120];
			end
			5'd16: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:128];
			end
			5'd17: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:136];
			end
			5'd18: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:144];
			end
			5'd19: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:152];
			end
			5'd20: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:160];
			end
			5'd21: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:168];
			end
			5'd22: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:176];
			end
			5'd23: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:184];
			end
			5'd24: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:192];
			end
			5'd25: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:200];
			end
			5'd26: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:208];
			end
			5'd27: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:216];
			end
			5'd28: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:224];
			end
			5'd29: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:232];
			end
			5'd30: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:240];
			end
			5'd31: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:248];
			end
			6'd32: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:256];
			end
			6'd33: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:264];
			end
			6'd34: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:272];
			end
			6'd35: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:280];
			end
			6'd36: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:288];
			end
			6'd37: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:296];
			end
			6'd38: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:304];
			end
			6'd39: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:312];
			end
			6'd40: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:320];
			end
			6'd41: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:328];
			end
			6'd42: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:336];
			end
			6'd43: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:344];
			end
			6'd44: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:352];
			end
			6'd45: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:360];
			end
			6'd46: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:368];
			end
			6'd47: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:376];
			end
			6'd48: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:384];
			end
			6'd49: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:392];
			end
			6'd50: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:400];
			end
			6'd51: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:408];
			end
			6'd52: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:416];
			end
			6'd53: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:424];
			end
			6'd54: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:432];
			end
			6'd55: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:440];
			end
			6'd56: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:448];
			end
			6'd57: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:456];
			end
			6'd58: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:464];
			end
			6'd59: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:472];
			end
			6'd60: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:480];
			end
			6'd61: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:488];
			end
			6'd62: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:496];
			end
			6'd63: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:504];
			end
			7'd64: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:512];
			end
			7'd65: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:520];
			end
			7'd66: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:528];
			end
			7'd67: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:536];
			end
			7'd68: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:544];
			end
			7'd69: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:552];
			end
			7'd70: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:560];
			end
			7'd71: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:568];
			end
			7'd72: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:576];
			end
			7'd73: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:584];
			end
			7'd74: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:592];
			end
			7'd75: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:600];
			end
			7'd76: begin
				monroe_ionphoton_dma_rawslicer_buf <= monroe_ionphoton_dma_rawslicer_buf[735:608];
			end
		endcase
	end
	clockdomainsrenamer_resetinserter_state <= clockdomainsrenamer_resetinserter_next_state;
	if (monroe_ionphoton_dma_reset) begin
		monroe_ionphoton_dma_rawslicer_buf <= 736'd0;
		monroe_ionphoton_dma_rawslicer_level <= 7'd0;
		clockdomainsrenamer_resetinserter_state <= 2'd0;
	end
	clockdomainsrenamer_recordconverter_state <= clockdomainsrenamer_recordconverter_next_state;
	if (monroe_ionphoton_dma_time_offset_source_ack) begin
		monroe_ionphoton_dma_time_offset_source_stb <= 1'd0;
	end
	if ((~monroe_ionphoton_dma_time_offset_source_stb)) begin
		monroe_ionphoton_dma_time_offset_source_payload_length <= monroe_ionphoton_dma_time_offset_sink_payload_length;
		monroe_ionphoton_dma_time_offset_source_payload_channel <= monroe_ionphoton_dma_time_offset_sink_payload_channel;
		monroe_ionphoton_dma_time_offset_source_payload_address <= monroe_ionphoton_dma_time_offset_sink_payload_address;
		monroe_ionphoton_dma_time_offset_source_payload_data <= monroe_ionphoton_dma_time_offset_sink_payload_data;
		monroe_ionphoton_dma_time_offset_source_payload_timestamp <= (monroe_ionphoton_dma_time_offset_sink_payload_timestamp + monroe_ionphoton_dma_time_offset_storage);
		monroe_ionphoton_dma_time_offset_source_eop <= monroe_ionphoton_dma_time_offset_sink_eop;
		monroe_ionphoton_dma_time_offset_source_stb <= monroe_ionphoton_dma_time_offset_sink_stb;
	end
	if (monroe_ionphoton_dma_cri_master_underflow_trigger) begin
		monroe_ionphoton_dma_cri_master_error_w <= 1'd1;
		monroe_ionphoton_dma_cri_master_error_channel_status <= monroe_ionphoton_dma_cri_master_sink_payload_channel;
		monroe_ionphoton_dma_cri_master_error_timestamp_status <= monroe_ionphoton_dma_cri_master_sink_payload_timestamp;
		monroe_ionphoton_dma_cri_master_error_address_status <= monroe_ionphoton_dma_cri_master_sink_payload_address;
	end
	if (monroe_ionphoton_dma_cri_master_link_error_trigger) begin
		monroe_ionphoton_dma_cri_master_error_w <= 2'd2;
		monroe_ionphoton_dma_cri_master_error_channel_status <= monroe_ionphoton_dma_cri_master_sink_payload_channel;
		monroe_ionphoton_dma_cri_master_error_timestamp_status <= monroe_ionphoton_dma_cri_master_sink_payload_timestamp;
		monroe_ionphoton_dma_cri_master_error_address_status <= monroe_ionphoton_dma_cri_master_sink_payload_address;
	end
	if (monroe_ionphoton_dma_cri_master_error_re) begin
		monroe_ionphoton_dma_cri_master_error_w <= 1'd0;
	end
	clockdomainsrenamer_crimaster_state <= clockdomainsrenamer_crimaster_next_state;
	clockdomainsrenamer_fsm_state <= clockdomainsrenamer_fsm_next_state;
	if (sys_kernel_rst) begin
		monroe_ionphoton_dma_dma_sink_stb <= 1'd0;
		monroe_ionphoton_dma_dma_sink_eop <= 1'd0;
		monroe_ionphoton_dma_dma_sink_payload_address <= 30'd0;
		monroe_ionphoton_dma_dma_source_eop <= 1'd0;
		monroe_ionphoton_dma_dma_source_payload_data <= 128'd0;
		monroe_ionphoton_dma_dma_data_reg_loaded <= 1'd0;
		monroe_ionphoton_dma_dma_enable_r <= 1'd0;
		monroe_ionphoton_dma_rawslicer_buf <= 736'd0;
		monroe_ionphoton_dma_rawslicer_level <= 7'd0;
		monroe_ionphoton_dma_time_offset_source_stb <= 1'd0;
		monroe_ionphoton_dma_time_offset_source_eop <= 1'd0;
		monroe_ionphoton_dma_time_offset_source_payload_length <= 8'd0;
		monroe_ionphoton_dma_time_offset_source_payload_channel <= 24'd0;
		monroe_ionphoton_dma_time_offset_source_payload_timestamp <= 64'd0;
		monroe_ionphoton_dma_time_offset_source_payload_address <= 8'd0;
		monroe_ionphoton_dma_time_offset_source_payload_data <= 512'd0;
		monroe_ionphoton_dma_cri_master_error_w <= 2'd0;
		monroe_ionphoton_dma_cri_master_error_channel_status <= 24'd0;
		monroe_ionphoton_dma_cri_master_error_timestamp_status <= 64'd0;
		monroe_ionphoton_dma_cri_master_error_address_status <= 16'd0;
		clockdomainsrenamer_resetinserter_state <= 2'd0;
		clockdomainsrenamer_recordconverter_state <= 2'd0;
		clockdomainsrenamer_crimaster_state <= 3'd0;
		clockdomainsrenamer_fsm_state <= 3'd0;
	end
end

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(23'd4194304)
) mor1kx (
	.clk(sys_clk),
	.dwbm_ack_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_ack),
	.dwbm_dat_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_r),
	.dwbm_err_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_interrupt),
	.iwbm_ack_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_ack),
	.iwbm_dat_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_r),
	.iwbm_err_i(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_rst),
	.dwbm_adr_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_d_adr_o),
	.dwbm_bte_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_bte),
	.dwbm_cti_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cti),
	.dwbm_cyc_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_cyc),
	.dwbm_dat_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_dat_w),
	.dwbm_sel_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_sel),
	.dwbm_stb_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_stb),
	.dwbm_we_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_dbus_we),
	.iwbm_adr_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_i_adr_o),
	.iwbm_bte_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_bte),
	.iwbm_cti_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cti),
	.iwbm_cyc_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_cyc),
	.iwbm_dat_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_dat_w),
	.iwbm_sel_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_sel),
	.iwbm_stb_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_stb),
	.iwbm_we_o(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ibus_we)
);

reg [31:0] mem[0:1023];
reg [9:0] memadr;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[0])
		mem[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr][7:0] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w[7:0];
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[1])
		mem[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr][15:8] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w[15:8];
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[2])
		mem[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr][23:16] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w[23:16];
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_we[3])
		mem[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr][31:24] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_w[31:24];
	memadr <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_sram_dat_r = mem[memadr];

reg [8:0] storage[0:15];
reg [8:0] memdat;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_we)
		storage[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_wrport_dat_r = memdat;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_dat_r = storage[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_tx_fifo_rdport_adr];

reg [8:0] storage_1[0:15];
reg [8:0] memdat_1;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_we)
		storage_1[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_dat_w;
	memdat_1 <= storage_1[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_wrport_dat_r = memdat_1;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_dat_r = storage_1[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_uart_rx_fifo_rdport_adr];

IBUFDS_GTE2 IBUFDS_GTE2(
	.CEB(1'd0),
	.I(clk125_gtp_p),
	.IB(clk125_gtp_n),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_buf),
	.ODIV2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_div2)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(14.5),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(8.0),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(90.0),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE (
	.CLKFBIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_fb),
	.CLKIN1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_div2),
	.CLKFBOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_fb),
	.CLKOUT0(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys),
	.CLKOUT1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x),
	.CLKOUT2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x_dqs),
	.LOCKED(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_locked)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE(3'd5),
	.CLKOUT0_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1)
) PLLE2_BASE (
	.CLKFBIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_fb),
	.CLKIN1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_div2),
	.CLKFBOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_fb),
	.CLKOUT0(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_clk200),
	.LOCKED(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_locked)
);

BUFG BUFG(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_2(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_mmcm_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

BUFG BUFG_3(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_pll_clk200),
	.O(clk200_clk)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg),
	.Q(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_meta),
	.PRE(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg),
	.Q(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_unbuf)
);

BUFG BUFG_4(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_asyncresetsynchronizerbufg_rst_unbuf),
	.O(sys_rst)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ic_reset)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[0]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[0]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[0]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[0]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[0]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[0]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[1]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[1]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[1]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[1]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[1]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[1]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[1]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[2]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[2]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[2]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[2]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[2]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[2]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[2]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[3]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[3]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[3]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[3]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[3]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[3]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[3]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[4]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[4]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[4]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[4]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[4]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[4]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[4]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[5]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[5]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[5]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[5]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[5]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[5]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[5]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[6]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[6]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[6]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[6]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[6]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[6]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[6]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[7]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[7]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[7]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[7]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[7]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[7]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[7]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[8]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[8]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[8]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[8]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[8]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[8]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[8]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[9]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[9]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[9]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[9]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[9]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[9]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[9]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[10]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[10]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[10]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[10]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[10]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[10]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[10]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[11]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[11]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[11]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[11]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[11]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[11]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[11]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[12]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[12]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[12]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[12]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[12]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[12]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[12]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[13]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[13]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[13]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[13]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[13]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[13]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[13]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[14]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_address[14]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[14]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_address[14]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[14]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_address[14]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[14]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[0]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[0]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[0]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[0]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[0]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[0]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[1]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[1]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[1]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[1]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[1]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[1]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[1]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[2]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_bank[2]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[2]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_bank[2]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[2]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_bank[2]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[2]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_ras_n),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_ras_n),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_ras_n),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_ras_n),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_ras_n),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_ras_n),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_ras_n),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cas_n),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cas_n),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cas_n),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cas_n),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cas_n),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cas_n),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cas_n),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_we_n),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_we_n),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_we_n),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_we_n),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_we_n),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_we_n),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_we_n),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cke),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_cke),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cke),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_cke),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cke),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_cke),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cke),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_odt),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_odt),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_odt),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_odt),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_odt),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_odt),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_odt),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_reset_n),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_reset_n),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_reset_n),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_reset_n),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_reset_n),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_reset_n),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_reset_n),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[1]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[2]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[3]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[4]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[5]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[6]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs0),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs0),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[1]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[2]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[3]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[4]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[5]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[6]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs1),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs1),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[0]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[16]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[0]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[16]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[0]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[16]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[0]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o0),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[16]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[0]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[16]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[0]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[16]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[0]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[16]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o0),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[1]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[17]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[1]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[17]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[1]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[17]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[1]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o1),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[17]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[1]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[17]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[1]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[17]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[1]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[17]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[1])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o1),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[2]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[18]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[2]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[18]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[2]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[18]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[2]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o2),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[18]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[2]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[18]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[2]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[18]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[2]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[18]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[2])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o2),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[3]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[19]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[3]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[19]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[3]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[19]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[3]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o3),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[19]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[3]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[19]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[3]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[19]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[3]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[19]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[3])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o3),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[4]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[20]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[4]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[20]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[4]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[20]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[4]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o4),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[20]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[4]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[20]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[4]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[20]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[4]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[20]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[4])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o4),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[5]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[21]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[5]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[21]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[5]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[21]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[5]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o5),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[21]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[5]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[21]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[5]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[21]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[5]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[21]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[5])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o5),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[6]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[22]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[6]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[22]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[6]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[22]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[6]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o6),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[22]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[6]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[22]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[6]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[22]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[6]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[22]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[6])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o6),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[7]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[23]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[7]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[23]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[7]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[23]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[7]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o7),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[23]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[7]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[23]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[7]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[23]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[7]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[23]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[7])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[0] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o7),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[8]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[24]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[8]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[24]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[8]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[24]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[8]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o8),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[24]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[8]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[24]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[8]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[24]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[8]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[24]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[8])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o8),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[9]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[25]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[9]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[25]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[9]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[25]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[9]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o9),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[25]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[9]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[25]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[9]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[25]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[9]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[25]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[9])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o9),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[10]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[26]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[10]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[26]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[10]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[26]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[10]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o10),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[26]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[10]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[26]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[10]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[26]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[10]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[26]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[10])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o10),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[11]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[27]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[11]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[27]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[11]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[27]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[11]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o11),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[27]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[11]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[27]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[11]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[27]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[11]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[27]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[11])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o11),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[12]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[28]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[12]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[28]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[12]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[28]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[12]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o12),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[28]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[12]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[28]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[12]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[28]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[12]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[28]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[12])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o12),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[13]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[29]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[13]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[29]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[13]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[29]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[13]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o13),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[29]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[13]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[29]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[13]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[29]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[13]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[29]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[13])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o13),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[14]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[30]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[14]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[30]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[14]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[30]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[14]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o14),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[30]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[14]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[30]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[14]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[30]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[14]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[30]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[14])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o14),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[15]),
	.D2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_wrdata[31]),
	.D3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[15]),
	.D4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_wrdata[31]),
	.D5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[15]),
	.D6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_wrdata[31]),
	.D7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[15]),
	.D8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o15),
	.TQ(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re))),
	.Q1(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[31]),
	.Q2(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p3_rddata[15]),
	.Q3(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[31]),
	.Q4(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p2_rddata[15]),
	.Q5(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[31]),
	.Q6(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p1_rddata[15]),
	.Q7(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[31]),
	.Q8(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dfi_p0_rddata[15])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_storage[1] & monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_o15),
	.T(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_ddrphy_dq_i_nodelay15)
);

reg [19:0] tag_mem[0:8191];
reg [12:0] memadr_1;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_we)
		tag_mem[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_w;
	memadr_1 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_tag_port_dat_r = tag_mem[memadr_1];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

assign spiflash2x_dq = monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_oe ? monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_o : 2'bz;
assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_spiflash_i0 = spiflash2x_dq;

GTPE2_COMMON #(
	.PLL0_FBDIV(3'd4),
	.PLL0_FBDIV_45(3'd5),
	.PLL0_REFCLK_DIV(1'd1)
) GTPE2_COMMON (
	.BGBYPASSB(1'd1),
	.BGMONITORENB(1'd1),
	.BGPDB(1'd1),
	.BGRCALOVRD(5'd31),
	.GTREFCLK0(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_clk125_buf),
	.GTREFCLK1(1'd0),
	.PLL0LOCKEN(1'd1),
	.PLL0PD(1'd0),
	.PLL0REFCLKSEL(1'd1),
	.PLL0RESET(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_reset),
	.PLL1PD(1'd1),
	.RCALENB(1'd1),
	.PLL0LOCK(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_lock),
	.PLL0OUTCLK(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_clk),
	.PLL0OUTREFCLK(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_refclk)
);

GTPE2_CHANNEL #(
	.ACJTAG_DEBUG_MODE(1'd0),
	.ACJTAG_MODE(1'd0),
	.ACJTAG_RESET(1'd0),
	.ADAPT_CFG0(1'd0),
	.ALIGN_COMMA_DOUBLE("FALSE"),
	.ALIGN_COMMA_ENABLE(10'd1023),
	.ALIGN_COMMA_WORD(1'd1),
	.ALIGN_MCOMMA_DET("TRUE"),
	.ALIGN_MCOMMA_VALUE(10'd643),
	.ALIGN_PCOMMA_DET("TRUE"),
	.ALIGN_PCOMMA_VALUE(9'd380),
	.CBCC_DATA_SOURCE_SEL("ENCODED"),
	.CFOK_CFG(43'd5016522067584),
	.CFOK_CFG2(6'd32),
	.CFOK_CFG3(6'd32),
	.CFOK_CFG4(1'd0),
	.CFOK_CFG5(1'd0),
	.CFOK_CFG6(1'd0),
	.CHAN_BOND_KEEP_ALIGN("FALSE"),
	.CHAN_BOND_MAX_SKEW(1'd1),
	.CHAN_BOND_SEQ_1_1(1'd0),
	.CHAN_BOND_SEQ_1_2(1'd0),
	.CHAN_BOND_SEQ_1_3(1'd0),
	.CHAN_BOND_SEQ_1_4(1'd0),
	.CHAN_BOND_SEQ_1_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_1(1'd0),
	.CHAN_BOND_SEQ_2_2(1'd0),
	.CHAN_BOND_SEQ_2_3(1'd0),
	.CHAN_BOND_SEQ_2_4(1'd0),
	.CHAN_BOND_SEQ_2_ENABLE(4'd15),
	.CHAN_BOND_SEQ_2_USE("FALSE"),
	.CHAN_BOND_SEQ_LEN(1'd1),
	.CLK_COMMON_SWING(1'd0),
	.CLK_CORRECT_USE("FALSE"),
	.CLK_COR_KEEP_IDLE("FALSE"),
	.CLK_COR_MAX_LAT(4'd9),
	.CLK_COR_MIN_LAT(3'd7),
	.CLK_COR_PRECEDENCE("TRUE"),
	.CLK_COR_REPEAT_WAIT(1'd0),
	.CLK_COR_SEQ_1_1(9'd256),
	.CLK_COR_SEQ_1_2(1'd0),
	.CLK_COR_SEQ_1_3(1'd0),
	.CLK_COR_SEQ_1_4(1'd0),
	.CLK_COR_SEQ_1_ENABLE(4'd15),
	.CLK_COR_SEQ_2_1(9'd256),
	.CLK_COR_SEQ_2_2(1'd0),
	.CLK_COR_SEQ_2_3(1'd0),
	.CLK_COR_SEQ_2_4(1'd0),
	.CLK_COR_SEQ_2_ENABLE(4'd15),
	.CLK_COR_SEQ_2_USE("FALSE"),
	.CLK_COR_SEQ_LEN(1'd1),
	.DEC_MCOMMA_DETECT("FALSE"),
	.DEC_PCOMMA_DETECT("FALSE"),
	.DEC_VALID_COMMA_ONLY("FALSE"),
	.DMONITOR_CFG(12'd2560),
	.ES_CLK_PHASE_SEL(1'd0),
	.ES_CONTROL(1'd0),
	.ES_ERRDET_EN("FALSE"),
	.ES_EYE_SCAN_EN("FALSE"),
	.ES_HORZ_OFFSET(5'd16),
	.ES_PMA_CFG(1'd0),
	.ES_PRESCALE(1'd0),
	.ES_QUALIFIER(1'd0),
	.ES_QUAL_MASK(1'd0),
	.ES_SDATA_MASK(1'd0),
	.ES_VERT_OFFSET(1'd0),
	.FTS_DESKEW_SEQ_ENABLE(4'd15),
	.FTS_LANE_DESKEW_CFG(4'd15),
	.FTS_LANE_DESKEW_EN("FALSE"),
	.GEARBOX_MODE(1'd0),
	.LOOPBACK_CFG(1'd0),
	.OUTREFCLK_SEL_INV(2'd3),
	.PCS_PCIE_EN("FALSE"),
	.PCS_RSVD_ATTR(1'd0),
	.PD_TRANS_TIME_FROM_P2(6'd60),
	.PD_TRANS_TIME_NONE_P2(6'd60),
	.PD_TRANS_TIME_TO_P2(7'd100),
	.PMA_LOOPBACK_CFG(1'd0),
	.PMA_RSV(10'd819),
	.PMA_RSV2(14'd8256),
	.PMA_RSV3(1'd0),
	.PMA_RSV4(1'd0),
	.PMA_RSV5(1'd0),
	.PMA_RSV6(1'd0),
	.PMA_RSV7(1'd0),
	.RXBUFRESET_TIME(1'd1),
	.RXBUF_ADDR_MODE("FAST"),
	.RXBUF_EIDLE_HI_CNT(4'd8),
	.RXBUF_EIDLE_LO_CNT(1'd0),
	.RXBUF_EN("TRUE"),
	.RXBUF_RESET_ON_CB_CHANGE("TRUE"),
	.RXBUF_RESET_ON_COMMAALIGN("FALSE"),
	.RXBUF_RESET_ON_EIDLE("FALSE"),
	.RXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.RXBUF_THRESH_OVFLW(6'd61),
	.RXBUF_THRESH_OVRD("FALSE"),
	.RXBUF_THRESH_UNDFLW(3'd4),
	.RXCDRFREQRESET_TIME(1'd1),
	.RXCDRPHRESET_TIME(1'd1),
	.RXCDR_CFG(69'd314170556264376963088),
	.RXCDR_FR_RESET_ON_EIDLE(1'd0),
	.RXCDR_HOLD_DURING_EIDLE(1'd0),
	.RXCDR_LOCK_CFG(4'd9),
	.RXCDR_PH_RESET_ON_EIDLE(1'd0),
	.RXDLY_CFG(5'd31),
	.RXDLY_LCFG(6'd48),
	.RXDLY_TAP_CFG(1'd0),
	.RXGEARBOX_EN("FALSE"),
	.RXISCANRESET_TIME(1'd1),
	.RXLPMRESET_TIME(4'd15),
	.RXLPM_BIAS_STARTUP_DISABLE(1'd0),
	.RXLPM_CFG(3'd6),
	.RXLPM_CFG1(1'd0),
	.RXLPM_CM_CFG(1'd0),
	.RXLPM_GC_CFG(9'd482),
	.RXLPM_GC_CFG2(1'd1),
	.RXLPM_HF_CFG(10'd1008),
	.RXLPM_HF_CFG2(4'd10),
	.RXLPM_HF_CFG3(1'd0),
	.RXLPM_HOLD_DURING_EIDLE(1'd0),
	.RXLPM_INCM_CFG(1'd0),
	.RXLPM_IPCM_CFG(1'd1),
	.RXLPM_LF_CFG(10'd1008),
	.RXLPM_LF_CFG2(4'd10),
	.RXLPM_OSINT_CFG(3'd4),
	.RXOOB_CFG(3'd6),
	.RXOOB_CLK_CFG("PMA"),
	.RXOSCALRESET_TIME(2'd3),
	.RXOSCALRESET_TIMEOUT(1'd0),
	.RXOUT_DIV(3'd4),
	.RXPCSRESET_TIME(1'd1),
	.RXPHDLY_CFG(20'd540704),
	.RXPH_CFG(24'd12582914),
	.RXPH_MONITOR_SEL(1'd0),
	.RXPI_CFG0(1'd0),
	.RXPI_CFG1(1'd1),
	.RXPI_CFG2(1'd1),
	.RXPMARESET_TIME(2'd3),
	.RXPRBS_ERR_LOOPBACK(1'd0),
	.RXSLIDE_AUTO_WAIT(3'd7),
	.RXSLIDE_MODE("OFF"),
	.RXSYNC_MULTILANE(1'd0),
	.RXSYNC_OVRD(1'd0),
	.RXSYNC_SKIP_DA(1'd0),
	.RX_BIAS_CFG(12'd3891),
	.RX_BUFFER_CFG(1'd0),
	.RX_CLK25_DIV(3'd5),
	.RX_CLKMUX_EN(1'd1),
	.RX_CM_SEL(1'd1),
	.RX_CM_TRIM(1'd0),
	.RX_DATA_WIDTH(5'd20),
	.RX_DDI_SEL(1'd0),
	.RX_DEBUG_CFG(1'd0),
	.RX_DEFER_RESET_BUF_EN("TRUE"),
	.RX_DISPERR_SEQ_MATCH("FALSE"),
	.RX_OS_CFG(8'd128),
	.RX_SIG_VALID_DLY(4'd10),
	.RX_XCLK_SEL("RXREC"),
	.SAS_MAX_COM(7'd64),
	.SAS_MIN_COM(6'd36),
	.SATA_BURST_SEQ_LEN(3'd5),
	.SATA_BURST_VAL(3'd4),
	.SATA_EIDLE_VAL(3'd4),
	.SATA_MAX_BURST(4'd8),
	.SATA_MAX_INIT(5'd21),
	.SATA_MAX_WAKE(3'd7),
	.SATA_MIN_BURST(3'd4),
	.SATA_MIN_INIT(4'd12),
	.SATA_MIN_WAKE(3'd4),
	.SATA_PLL_CFG("VCO_3000MHZ"),
	.SHOW_REALIGN_COMMA("TRUE"),
	.SIM_RECEIVER_DETECT_PASS("TRUE"),
	.SIM_RESET_SPEEDUP("FALSE"),
	.SIM_TX_EIDLE_DRIVE_LEVEL("X"),
	.SIM_VERSION("2.0"),
	.TERM_RCAL_CFG(15'd16912),
	.TERM_RCAL_OVRD(1'd0),
	.TRANS_TIME_RATE(4'd14),
	.TST_RSV(1'd0),
	.TXBUF_EN("TRUE"),
	.TXBUF_RESET_ON_RATE_CHANGE("TRUE"),
	.TXDLY_CFG(5'd31),
	.TXDLY_LCFG(6'd48),
	.TXDLY_TAP_CFG(1'd0),
	.TXGEARBOX_EN("FALSE"),
	.TXOOB_CFG(1'd0),
	.TXOUT_DIV(3'd4),
	.TXPCSRESET_TIME(1'd1),
	.TXPHDLY_CFG(20'd540704),
	.TXPH_CFG(11'd1920),
	.TXPH_MONITOR_SEL(1'd0),
	.TXPI_CFG0(1'd0),
	.TXPI_CFG1(1'd0),
	.TXPI_CFG2(1'd0),
	.TXPI_CFG3(1'd0),
	.TXPI_CFG4(1'd0),
	.TXPI_CFG5(1'd0),
	.TXPI_GREY_SEL(1'd0),
	.TXPI_INVSTROBE_SEL(1'd0),
	.TXPI_PPMCLK_SEL("TXUSRCLK2"),
	.TXPI_PPM_CFG(1'd0),
	.TXPI_SYNFREQ_PPM(1'd1),
	.TXPMARESET_TIME(1'd1),
	.TXSYNC_MULTILANE(1'd0),
	.TXSYNC_OVRD(1'd0),
	.TXSYNC_SKIP_DA(1'd0),
	.TX_CLK25_DIV(3'd5),
	.TX_CLKMUX_EN(1'd1),
	.TX_DATA_WIDTH(5'd20),
	.TX_DEEMPH0(1'd0),
	.TX_DEEMPH1(1'd0),
	.TX_DRIVE_MODE("DIRECT"),
	.TX_EIDLE_ASSERT_DELAY(3'd6),
	.TX_EIDLE_DEASSERT_DELAY(3'd4),
	.TX_LOOPBACK_DRIVE_HIZ("FALSE"),
	.TX_MAINCURSOR_SEL(1'd0),
	.TX_MARGIN_FULL_0(7'd78),
	.TX_MARGIN_FULL_1(7'd73),
	.TX_MARGIN_FULL_2(7'd69),
	.TX_MARGIN_FULL_3(7'd66),
	.TX_MARGIN_FULL_4(7'd64),
	.TX_MARGIN_LOW_0(7'd70),
	.TX_MARGIN_LOW_1(7'd68),
	.TX_MARGIN_LOW_2(7'd66),
	.TX_MARGIN_LOW_3(7'd64),
	.TX_MARGIN_LOW_4(7'd64),
	.TX_PREDRIVER_MODE(1'd0),
	.TX_RXDETECT_CFG(13'd6194),
	.TX_RXDETECT_REF(3'd4),
	.TX_XCLK_SEL("TXOUT"),
	.UCODEER_CLR(1'd0),
	.USE_PCS_CLK_PHASE_SEL(1'd0)
) GTPE2_CHANNEL (
	.CFGRESET(1'd0),
	.CLKRSVD0(1'd0),
	.CLKRSVD1(1'd0),
	.DMONFIFORESET(1'd0),
	.DMONITORCLK(1'd0),
	.DRPADDR(monroe_ionphoton_monroe_ionphoton_drpaddr),
	.DRPCLK(sys_clk),
	.DRPDI(monroe_ionphoton_monroe_ionphoton_drpdi),
	.DRPEN(monroe_ionphoton_monroe_ionphoton_drpen),
	.DRPWE(monroe_ionphoton_monroe_ionphoton_drpwe),
	.EYESCANMODE(1'd0),
	.EYESCANRESET(1'd0),
	.EYESCANTRIGGER(1'd0),
	.GTPRXN(sfp_rxn),
	.GTPRXP(sfp_rxp),
	.GTRESETSEL(1'd0),
	.GTRSVD(1'd0),
	.GTRXRESET(monroe_ionphoton_monroe_ionphoton_rx_reset),
	.GTTXRESET(monroe_ionphoton_monroe_ionphoton_tx_reset),
	.LOOPBACK(1'd0),
	.PCSRSVDIN(1'd0),
	.PLL0CLK(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_clk),
	.PLL0REFCLK(monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_qpll_refclk),
	.PLL1CLK(1'd0),
	.PLL1REFCLK(1'd0),
	.PMARSVDIN0(1'd0),
	.PMARSVDIN1(1'd0),
	.PMARSVDIN2(1'd0),
	.PMARSVDIN3(1'd0),
	.PMARSVDIN4(1'd0),
	.RESETOVRD(1'd0),
	.RX8B10BEN(1'd0),
	.RXADAPTSELTEST(1'd0),
	.RXBUFRESET(1'd0),
	.RXCDRFREQRESET(1'd0),
	.RXCDRHOLD(1'd0),
	.RXCDROVRDEN(1'd0),
	.RXCDRRESET(1'd0),
	.RXCDRRESETRSV(1'd0),
	.RXCHBONDEN(1'd0),
	.RXCHBONDI(1'd0),
	.RXCHBONDLEVEL(1'd0),
	.RXCHBONDMASTER(1'd0),
	.RXCHBONDSLAVE(1'd0),
	.RXCOMMADETEN(1'd0),
	.RXDDIEN(1'd0),
	.RXDFEXYDEN(1'd0),
	.RXDLYBYPASS(1'd1),
	.RXDLYEN(1'd0),
	.RXDLYOVRDEN(1'd0),
	.RXDLYSRESET(1'd0),
	.RXELECIDLEMODE(2'd3),
	.RXGEARBOXSLIP(1'd0),
	.RXLPMHFHOLD(1'd0),
	.RXLPMHFOVRDEN(1'd0),
	.RXLPMLFHOLD(1'd0),
	.RXLPMLFOVRDEN(1'd0),
	.RXLPMOSINTNTRLEN(1'd0),
	.RXLPMRESET(1'd0),
	.RXMCOMMAALIGNEN(1'd0),
	.RXOOBRESET(1'd0),
	.RXOSCALRESET(1'd0),
	.RXOSHOLD(1'd0),
	.RXOSINTCFG(2'd2),
	.RXOSINTEN(1'd1),
	.RXOSINTHOLD(1'd0),
	.RXOSINTID0(1'd0),
	.RXOSINTNTRLEN(1'd0),
	.RXOSINTOVRDEN(1'd0),
	.RXOSINTPD(1'd0),
	.RXOSINTSTROBE(1'd0),
	.RXOSINTTESTOVRDEN(1'd0),
	.RXOSOVRDEN(1'd0),
	.RXOUTCLKSEL(2'd2),
	.RXPCOMMAALIGNEN(1'd0),
	.RXPCSRESET(1'd0),
	.RXPD(1'd0),
	.RXPHALIGN(1'd0),
	.RXPHALIGNEN(1'd0),
	.RXPHDLYPD(1'd0),
	.RXPHDLYRESET(1'd0),
	.RXPHOVRDEN(1'd0),
	.RXPMARESET(1'd0),
	.RXPOLARITY(1'd0),
	.RXPRBSCNTRESET(1'd0),
	.RXPRBSSEL(1'd0),
	.RXRATE(1'd0),
	.RXRATEMODE(1'd0),
	.RXSLIDE(1'd0),
	.RXSYNCALLIN(1'd0),
	.RXSYNCIN(1'd0),
	.RXSYNCMODE(1'd0),
	.RXSYSCLKSEL(1'd0),
	.RXUSERRDY(monroe_ionphoton_monroe_ionphoton_rx_mmcm_locked),
	.RXUSRCLK(eth_rx_half_clk),
	.RXUSRCLK2(eth_rx_half_clk),
	.SETERRSTATUS(1'd0),
	.SIGVALIDCLK(1'd0),
	.TSTIN(20'd1048575),
	.TX8B10BBYPASS(1'd0),
	.TX8B10BEN(1'd0),
	.TXBUFDIFFCTRL(3'd4),
	.TXCHARDISPMODE({monroe_ionphoton_monroe_ionphoton_tx_data0[19], monroe_ionphoton_monroe_ionphoton_tx_data0[9]}),
	.TXCHARDISPVAL({monroe_ionphoton_monroe_ionphoton_tx_data0[18], monroe_ionphoton_monroe_ionphoton_tx_data0[8]}),
	.TXCHARISK(1'd0),
	.TXCOMINIT(1'd0),
	.TXCOMSAS(1'd0),
	.TXCOMWAKE(1'd0),
	.TXDATA({monroe_ionphoton_monroe_ionphoton_tx_data0[17:10], monroe_ionphoton_monroe_ionphoton_tx_data0[7:0]}),
	.TXDEEMPH(1'd0),
	.TXDETECTRX(1'd0),
	.TXDIFFCTRL(4'd8),
	.TXDIFFPD(1'd0),
	.TXDLYBYPASS(1'd1),
	.TXDLYEN(1'd0),
	.TXDLYHOLD(1'd0),
	.TXDLYOVRDEN(1'd0),
	.TXDLYSRESET(1'd0),
	.TXDLYUPDOWN(1'd0),
	.TXELECIDLE(1'd0),
	.TXHEADER(1'd0),
	.TXINHIBIT(1'd0),
	.TXMAINCURSOR(1'd0),
	.TXMARGIN(1'd0),
	.TXOUTCLKSEL(2'd2),
	.TXPCSRESET(1'd0),
	.TXPD(1'd0),
	.TXPDELECIDLEMODE(1'd0),
	.TXPHALIGN(1'd0),
	.TXPHALIGNEN(1'd0),
	.TXPHDLYPD(1'd0),
	.TXPHDLYRESET(1'd0),
	.TXPHDLYTSTCLK(1'd0),
	.TXPHINIT(1'd0),
	.TXPHOVRDEN(1'd0),
	.TXPIPPMEN(1'd0),
	.TXPIPPMOVRDEN(1'd0),
	.TXPIPPMPD(1'd0),
	.TXPIPPMSEL(1'd1),
	.TXPIPPMSTEPSIZE(1'd0),
	.TXPISOPD(1'd0),
	.TXPMARESET(1'd0),
	.TXPOLARITY(1'd0),
	.TXPOSTCURSOR(1'd0),
	.TXPOSTCURSORINV(1'd0),
	.TXPRBSFORCEERR(1'd0),
	.TXPRBSSEL(1'd0),
	.TXPRECURSOR(1'd0),
	.TXPRECURSORINV(1'd0),
	.TXRATE(1'd0),
	.TXRATEMODE(1'd0),
	.TXSEQUENCE(1'd0),
	.TXSTARTSEQ(1'd0),
	.TXSWING(1'd0),
	.TXSYNCALLIN(1'd0),
	.TXSYNCIN(1'd0),
	.TXSYNCMODE(1'd0),
	.TXSYSCLKSEL(1'd0),
	.TXUSERRDY(monroe_ionphoton_monroe_ionphoton_tx_mmcm_locked),
	.TXUSRCLK(eth_tx_half_clk),
	.TXUSRCLK2(eth_tx_half_clk),
	.DRPDO(monroe_ionphoton_monroe_ionphoton_drpdo),
	.DRPRDY(monroe_ionphoton_monroe_ionphoton_drprdy),
	.GTPTXN(sfp_txn),
	.GTPTXP(sfp_txp),
	.RXCHARISK({monroe_ionphoton_monroe_ionphoton_rx_data0[18], monroe_ionphoton_monroe_ionphoton_rx_data0[8]}),
	.RXDATA({monroe_ionphoton_monroe_ionphoton_rx_data0[17:10], monroe_ionphoton_monroe_ionphoton_rx_data0[7:0]}),
	.RXDISPERR({monroe_ionphoton_monroe_ionphoton_rx_data0[19], monroe_ionphoton_monroe_ionphoton_rx_data0[9]}),
	.RXOUTCLK(monroe_ionphoton_monroe_ionphoton_rxoutclk),
	.RXPMARESETDONE(monroe_ionphoton_monroe_ionphoton_rx_pma_reset_done),
	.RXRESETDONE(monroe_ionphoton_monroe_ionphoton_rx_reset_done),
	.TXOUTCLK(monroe_ionphoton_monroe_ionphoton_txoutclk),
	.TXRESETDONE(monroe_ionphoton_monroe_ionphoton_tx_reset_done)
);

BUFH BUFH(
	.I(monroe_ionphoton_monroe_ionphoton_txoutclk),
	.O(monroe_ionphoton_monroe_ionphoton_txoutclk_rebuffer)
);

BUFG BUFG_5(
	.I(monroe_ionphoton_monroe_ionphoton_rxoutclk),
	.O(monroe_ionphoton_monroe_ionphoton_rxoutclk_rebuffer)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE_1 (
	.CLKFBIN(monroe_ionphoton_monroe_ionphoton_tx_mmcm_fb),
	.CLKIN1(monroe_ionphoton_monroe_ionphoton_txoutclk_rebuffer),
	.RST(monroe_ionphoton_monroe_ionphoton_tx_mmcm_reset),
	.CLKFBOUT(monroe_ionphoton_monroe_ionphoton_tx_mmcm_fb),
	.CLKOUT0(monroe_ionphoton_monroe_ionphoton_clk_tx_half_unbuf),
	.CLKOUT1(monroe_ionphoton_monroe_ionphoton_clk_tx_unbuf),
	.LOCKED(monroe_ionphoton_monroe_ionphoton_tx_mmcm_locked)
);

BUFH BUFH_1(
	.I(monroe_ionphoton_monroe_ionphoton_clk_tx_half_unbuf),
	.O(eth_tx_half_clk)
);

BUFH BUFH_2(
	.I(monroe_ionphoton_monroe_ionphoton_clk_tx_unbuf),
	.O(eth_tx_clk)
);

MMCME2_BASE #(
	.CLKFBOUT_MULT_F(5'd16),
	.CLKIN1_PERIOD(16.0),
	.CLKOUT0_DIVIDE_F(5'd16),
	.CLKOUT1_DIVIDE(4'd8),
	.DIVCLK_DIVIDE(1'd1)
) MMCME2_BASE_2 (
	.CLKFBIN(monroe_ionphoton_monroe_ionphoton_rx_mmcm_fb),
	.CLKIN1(monroe_ionphoton_monroe_ionphoton_rxoutclk_rebuffer),
	.RST(monroe_ionphoton_monroe_ionphoton_rx_mmcm_reset),
	.CLKFBOUT(monroe_ionphoton_monroe_ionphoton_rx_mmcm_fb),
	.CLKOUT0(monroe_ionphoton_monroe_ionphoton_clk_rx_half_unbuf),
	.CLKOUT1(monroe_ionphoton_monroe_ionphoton_clk_rx_unbuf),
	.LOCKED(monroe_ionphoton_monroe_ionphoton_rx_mmcm_locked)
);

BUFG BUFG_6(
	.I(monroe_ionphoton_monroe_ionphoton_clk_rx_half_unbuf),
	.O(eth_rx_half_clk)
);

BUFG BUFG_7(
	.I(monroe_ionphoton_monroe_ionphoton_clk_rx_unbuf),
	.O(eth_rx_clk)
);

reg [10:0] storage_2[0:4];
reg [10:0] memdat_2;
always @(posedge eth_rx_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_we)
		storage_2[monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_dat_w;
	memdat_2 <= storage_2[monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_adr];
end

always @(posedge eth_rx_clk) begin
end

assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_wrport_dat_r = memdat_2;
assign monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_dat_r = storage_2[monroe_ionphoton_monroe_ionphoton_crc32_checker_syncfifo_rdport_adr];

reg [40:0] storage_3[0:63];
reg [5:0] memadr_2;
reg [5:0] memadr_3;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_we)
		storage_3[monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_dat_w;
	memadr_2 <= monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memadr_3 <= monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_adr;
end

assign monroe_ionphoton_monroe_ionphoton_tx_cdc_wrport_dat_r = storage_3[memadr_2];
assign monroe_ionphoton_monroe_ionphoton_tx_cdc_rdport_dat_r = storage_3[memadr_3];

reg [40:0] storage_4[0:63];
reg [5:0] memadr_4;
reg [5:0] memadr_5;
always @(posedge eth_rx_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_we)
		storage_4[monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_dat_w;
	memadr_4 <= monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_5 <= monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_adr;
end

assign monroe_ionphoton_monroe_ionphoton_rx_cdc_wrport_dat_r = storage_4[memadr_4];
assign monroe_ionphoton_monroe_ionphoton_rx_cdc_rdport_dat_r = storage_4[memadr_5];

reg [34:0] storage_5[0:3];
reg [34:0] memdat_3;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_we)
		storage_5[monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_dat_w;
	memdat_3 <= storage_5[monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign monroe_ionphoton_monroe_ionphoton_writer_fifo_wrport_dat_r = memdat_3;
assign monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_dat_r = storage_5[monroe_ionphoton_monroe_ionphoton_writer_fifo_rdport_adr];

reg [31:0] mem_1[0:381];
reg [8:0] memadr_6;
reg [8:0] memadr_7;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_writer_memory0_we)
		mem_1[monroe_ionphoton_monroe_ionphoton_writer_memory0_adr] <= monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_w;
	memadr_6 <= monroe_ionphoton_monroe_ionphoton_writer_memory0_adr;
end

always @(posedge sys_clk) begin
	memadr_7 <= monroe_ionphoton_monroe_ionphoton_sram0_adr0;
end

assign monroe_ionphoton_monroe_ionphoton_writer_memory0_dat_r = mem_1[memadr_6];
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_r0 = mem_1[memadr_7];

reg [31:0] mem_2[0:381];
reg [8:0] memadr_8;
reg [8:0] memadr_9;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_writer_memory1_we)
		mem_2[monroe_ionphoton_monroe_ionphoton_writer_memory1_adr] <= monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_w;
	memadr_8 <= monroe_ionphoton_monroe_ionphoton_writer_memory1_adr;
end

always @(posedge sys_clk) begin
	memadr_9 <= monroe_ionphoton_monroe_ionphoton_sram1_adr0;
end

assign monroe_ionphoton_monroe_ionphoton_writer_memory1_dat_r = mem_2[memadr_8];
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_r0 = mem_2[memadr_9];

reg [31:0] mem_3[0:381];
reg [8:0] memadr_10;
reg [8:0] memadr_11;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_writer_memory2_we)
		mem_3[monroe_ionphoton_monroe_ionphoton_writer_memory2_adr] <= monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_w;
	memadr_10 <= monroe_ionphoton_monroe_ionphoton_writer_memory2_adr;
end

always @(posedge sys_clk) begin
	memadr_11 <= monroe_ionphoton_monroe_ionphoton_sram2_adr0;
end

assign monroe_ionphoton_monroe_ionphoton_writer_memory2_dat_r = mem_3[memadr_10];
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_r0 = mem_3[memadr_11];

reg [31:0] mem_4[0:381];
reg [8:0] memadr_12;
reg [8:0] memadr_13;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_writer_memory3_we)
		mem_4[monroe_ionphoton_monroe_ionphoton_writer_memory3_adr] <= monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_w;
	memadr_12 <= monroe_ionphoton_monroe_ionphoton_writer_memory3_adr;
end

always @(posedge sys_clk) begin
	memadr_13 <= monroe_ionphoton_monroe_ionphoton_sram3_adr0;
end

assign monroe_ionphoton_monroe_ionphoton_writer_memory3_dat_r = mem_4[memadr_12];
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_r0 = mem_4[memadr_13];

reg [13:0] storage_6[0:3];
reg [13:0] memdat_4;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_we)
		storage_6[monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr] <= monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_dat_w;
	memdat_4 <= storage_6[monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign monroe_ionphoton_monroe_ionphoton_reader_fifo_wrport_dat_r = memdat_4;
assign monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_dat_r = storage_6[monroe_ionphoton_monroe_ionphoton_reader_fifo_rdport_adr];

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(31'd1082130432)
) mor1kx_1 (
	.clk(sys_kernel_clk),
	.dwbm_ack_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_ack),
	.dwbm_dat_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_r),
	.dwbm_err_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_interrupt),
	.iwbm_ack_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_ack),
	.iwbm_dat_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_r),
	.iwbm_err_i(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_kernel_rst),
	.dwbm_adr_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_d_adr_o),
	.dwbm_bte_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_bte),
	.dwbm_cti_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cti),
	.dwbm_cyc_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_cyc),
	.dwbm_dat_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_dat_w),
	.dwbm_sel_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_sel),
	.dwbm_stb_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_stb),
	.dwbm_we_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_dbus_we),
	.iwbm_adr_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_i_adr_o),
	.iwbm_bte_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_bte),
	.iwbm_cti_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cti),
	.iwbm_cyc_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_cyc),
	.iwbm_dat_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_dat_w),
	.iwbm_sel_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_sel),
	.iwbm_stb_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_stb),
	.iwbm_we_o(monroe_ionphoton_monroe_ionphoton_kernel_cpu_ibus_we)
);

reg [7:0] mem_5[0:37];
reg [5:0] memadr_14;
always @(posedge sys_clk) begin
	memadr_14 <= monroe_ionphoton_add_identifier_adr;
end

assign monroe_ionphoton_add_identifier_dat_r = mem_5[memadr_14];

initial begin
	$readmemh("mem_5.init", mem_5);
end

assign i2c_scl = monroe_ionphoton_i2c_tstriple0_oe ? monroe_ionphoton_i2c_tstriple0_o : 1'bz;
assign monroe_ionphoton_i2c_tstriple0_i = i2c_scl;

assign i2c_sda = monroe_ionphoton_i2c_tstriple1_oe ? monroe_ionphoton_i2c_tstriple1_o : 1'bz;
assign monroe_ionphoton_i2c_tstriple1_i = i2c_sda;

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_16 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(inout_8x0_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(inout_8x0_serdes_i1[7]),
	.Q2(inout_8x0_serdes_i1[6]),
	.Q3(inout_8x0_serdes_i1[5]),
	.Q4(inout_8x0_serdes_i1[4]),
	.Q5(inout_8x0_serdes_i1[3]),
	.Q6(inout_8x0_serdes_i1[2]),
	.Q7(inout_8x0_serdes_i1[1]),
	.Q8(inout_8x0_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(inout_8x0_serdes_o1[0]),
	.D2(inout_8x0_serdes_o1[1]),
	.D3(inout_8x0_serdes_o1[2]),
	.D4(inout_8x0_serdes_o1[3]),
	.D5(inout_8x0_serdes_o1[4]),
	.D6(inout_8x0_serdes_o1[5]),
	.D7(inout_8x0_serdes_o1[6]),
	.D8(inout_8x0_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(inout_8x0_serdes_t_in),
	.TCE(1'd1),
	.OQ(inout_8x0_serdes_pad_o1),
	.TQ(inout_8x0_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE (
	.I(inout_8x0_serdes_pad_o0),
	.IBUFDISABLE((~inout_8x0_serdes_t_out)),
	.INTERMDISABLE((~inout_8x0_serdes_t_out)),
	.T(inout_8x0_serdes_t_out),
	.IO(dio0_p),
	.IOB(dio0_n),
	.O(inout_8x0_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_17 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(inout_8x1_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(inout_8x1_serdes_i1[7]),
	.Q2(inout_8x1_serdes_i1[6]),
	.Q3(inout_8x1_serdes_i1[5]),
	.Q4(inout_8x1_serdes_i1[4]),
	.Q5(inout_8x1_serdes_i1[3]),
	.Q6(inout_8x1_serdes_i1[2]),
	.Q7(inout_8x1_serdes_i1[1]),
	.Q8(inout_8x1_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(inout_8x1_serdes_o1[0]),
	.D2(inout_8x1_serdes_o1[1]),
	.D3(inout_8x1_serdes_o1[2]),
	.D4(inout_8x1_serdes_o1[3]),
	.D5(inout_8x1_serdes_o1[4]),
	.D6(inout_8x1_serdes_o1[5]),
	.D7(inout_8x1_serdes_o1[6]),
	.D8(inout_8x1_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(inout_8x1_serdes_t_in),
	.TCE(1'd1),
	.OQ(inout_8x1_serdes_pad_o1),
	.TQ(inout_8x1_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_1 (
	.I(inout_8x1_serdes_pad_o0),
	.IBUFDISABLE((~inout_8x1_serdes_t_out)),
	.INTERMDISABLE((~inout_8x1_serdes_t_out)),
	.T(inout_8x1_serdes_t_out),
	.IO(dio0_p_1),
	.IOB(dio0_n_1),
	.O(inout_8x1_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_18 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(inout_8x2_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(inout_8x2_serdes_i1[7]),
	.Q2(inout_8x2_serdes_i1[6]),
	.Q3(inout_8x2_serdes_i1[5]),
	.Q4(inout_8x2_serdes_i1[4]),
	.Q5(inout_8x2_serdes_i1[3]),
	.Q6(inout_8x2_serdes_i1[2]),
	.Q7(inout_8x2_serdes_i1[1]),
	.Q8(inout_8x2_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(inout_8x2_serdes_o1[0]),
	.D2(inout_8x2_serdes_o1[1]),
	.D3(inout_8x2_serdes_o1[2]),
	.D4(inout_8x2_serdes_o1[3]),
	.D5(inout_8x2_serdes_o1[4]),
	.D6(inout_8x2_serdes_o1[5]),
	.D7(inout_8x2_serdes_o1[6]),
	.D8(inout_8x2_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(inout_8x2_serdes_t_in),
	.TCE(1'd1),
	.OQ(inout_8x2_serdes_pad_o1),
	.TQ(inout_8x2_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_2 (
	.I(inout_8x2_serdes_pad_o0),
	.IBUFDISABLE((~inout_8x2_serdes_t_out)),
	.INTERMDISABLE((~inout_8x2_serdes_t_out)),
	.T(inout_8x2_serdes_t_out),
	.IO(dio0_p_2),
	.IOB(dio0_n_2),
	.O(inout_8x2_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_19 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(inout_8x3_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(inout_8x3_serdes_i1[7]),
	.Q2(inout_8x3_serdes_i1[6]),
	.Q3(inout_8x3_serdes_i1[5]),
	.Q4(inout_8x3_serdes_i1[4]),
	.Q5(inout_8x3_serdes_i1[3]),
	.Q6(inout_8x3_serdes_i1[2]),
	.Q7(inout_8x3_serdes_i1[1]),
	.Q8(inout_8x3_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(inout_8x3_serdes_o1[0]),
	.D2(inout_8x3_serdes_o1[1]),
	.D3(inout_8x3_serdes_o1[2]),
	.D4(inout_8x3_serdes_o1[3]),
	.D5(inout_8x3_serdes_o1[4]),
	.D6(inout_8x3_serdes_o1[5]),
	.D7(inout_8x3_serdes_o1[6]),
	.D8(inout_8x3_serdes_o1[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(inout_8x3_serdes_t_in),
	.TCE(1'd1),
	.OQ(inout_8x3_serdes_pad_o1),
	.TQ(inout_8x3_serdes_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_3 (
	.I(inout_8x3_serdes_pad_o0),
	.IBUFDISABLE((~inout_8x3_serdes_t_out)),
	.INTERMDISABLE((~inout_8x3_serdes_t_out)),
	.T(inout_8x3_serdes_t_out),
	.IO(dio0_p_3),
	.IOB(dio0_n_3),
	.O(inout_8x3_serdes_pad_i0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x0_o[0]),
	.D2(output_8x0_o[1]),
	.D3(output_8x0_o[2]),
	.D4(output_8x0_o[3]),
	.D5(output_8x0_o[4]),
	.D6(output_8x0_o[5]),
	.D7(output_8x0_o[6]),
	.D8(output_8x0_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x0_t_in),
	.TCE(1'd1),
	.OQ(output_8x0_pad_o),
	.TQ(output_8x0_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_4 (
	.I(output_8x0_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x0_t_out),
	.IO(dio0_p_4),
	.IOB(dio0_n_4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x1_o[0]),
	.D2(output_8x1_o[1]),
	.D3(output_8x1_o[2]),
	.D4(output_8x1_o[3]),
	.D5(output_8x1_o[4]),
	.D6(output_8x1_o[5]),
	.D7(output_8x1_o[6]),
	.D8(output_8x1_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x1_t_in),
	.TCE(1'd1),
	.OQ(output_8x1_pad_o),
	.TQ(output_8x1_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_5 (
	.I(output_8x1_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x1_t_out),
	.IO(dio0_p_5),
	.IOB(dio0_n_5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x2_o[0]),
	.D2(output_8x2_o[1]),
	.D3(output_8x2_o[2]),
	.D4(output_8x2_o[3]),
	.D5(output_8x2_o[4]),
	.D6(output_8x2_o[5]),
	.D7(output_8x2_o[6]),
	.D8(output_8x2_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x2_t_in),
	.TCE(1'd1),
	.OQ(output_8x2_pad_o),
	.TQ(output_8x2_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_6 (
	.I(output_8x2_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x2_t_out),
	.IO(dio0_p_6),
	.IOB(dio0_n_6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x3_o[0]),
	.D2(output_8x3_o[1]),
	.D3(output_8x3_o[2]),
	.D4(output_8x3_o[3]),
	.D5(output_8x3_o[4]),
	.D6(output_8x3_o[5]),
	.D7(output_8x3_o[6]),
	.D8(output_8x3_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x3_t_in),
	.TCE(1'd1),
	.OQ(output_8x3_pad_o),
	.TQ(output_8x3_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_7 (
	.I(output_8x3_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x3_t_out),
	.IO(dio0_p_7),
	.IOB(dio0_n_7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_53 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x4_o[0]),
	.D2(output_8x4_o[1]),
	.D3(output_8x4_o[2]),
	.D4(output_8x4_o[3]),
	.D5(output_8x4_o[4]),
	.D6(output_8x4_o[5]),
	.D7(output_8x4_o[6]),
	.D8(output_8x4_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x4_t_in),
	.TCE(1'd1),
	.OQ(output_8x4_pad_o),
	.TQ(output_8x4_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_8 (
	.I(output_8x4_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x4_t_out),
	.IO(dio1_p),
	.IOB(dio1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_54 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x5_o[0]),
	.D2(output_8x5_o[1]),
	.D3(output_8x5_o[2]),
	.D4(output_8x5_o[3]),
	.D5(output_8x5_o[4]),
	.D6(output_8x5_o[5]),
	.D7(output_8x5_o[6]),
	.D8(output_8x5_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x5_t_in),
	.TCE(1'd1),
	.OQ(output_8x5_pad_o),
	.TQ(output_8x5_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_9 (
	.I(output_8x5_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x5_t_out),
	.IO(dio1_p_1),
	.IOB(dio1_n_1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_55 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x6_o[0]),
	.D2(output_8x6_o[1]),
	.D3(output_8x6_o[2]),
	.D4(output_8x6_o[3]),
	.D5(output_8x6_o[4]),
	.D6(output_8x6_o[5]),
	.D7(output_8x6_o[6]),
	.D8(output_8x6_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x6_t_in),
	.TCE(1'd1),
	.OQ(output_8x6_pad_o),
	.TQ(output_8x6_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_10 (
	.I(output_8x6_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x6_t_out),
	.IO(dio1_p_2),
	.IOB(dio1_n_2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_56 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x7_o[0]),
	.D2(output_8x7_o[1]),
	.D3(output_8x7_o[2]),
	.D4(output_8x7_o[3]),
	.D5(output_8x7_o[4]),
	.D6(output_8x7_o[5]),
	.D7(output_8x7_o[6]),
	.D8(output_8x7_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x7_t_in),
	.TCE(1'd1),
	.OQ(output_8x7_pad_o),
	.TQ(output_8x7_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_11 (
	.I(output_8x7_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x7_t_out),
	.IO(dio1_p_3),
	.IOB(dio1_n_3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_57 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x8_o[0]),
	.D2(output_8x8_o[1]),
	.D3(output_8x8_o[2]),
	.D4(output_8x8_o[3]),
	.D5(output_8x8_o[4]),
	.D6(output_8x8_o[5]),
	.D7(output_8x8_o[6]),
	.D8(output_8x8_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x8_t_in),
	.TCE(1'd1),
	.OQ(output_8x8_pad_o),
	.TQ(output_8x8_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_12 (
	.I(output_8x8_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x8_t_out),
	.IO(dio1_p_4),
	.IOB(dio1_n_4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_58 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x9_o[0]),
	.D2(output_8x9_o[1]),
	.D3(output_8x9_o[2]),
	.D4(output_8x9_o[3]),
	.D5(output_8x9_o[4]),
	.D6(output_8x9_o[5]),
	.D7(output_8x9_o[6]),
	.D8(output_8x9_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x9_t_in),
	.TCE(1'd1),
	.OQ(output_8x9_pad_o),
	.TQ(output_8x9_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_13 (
	.I(output_8x9_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x9_t_out),
	.IO(dio1_p_5),
	.IOB(dio1_n_5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_59 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x10_o[0]),
	.D2(output_8x10_o[1]),
	.D3(output_8x10_o[2]),
	.D4(output_8x10_o[3]),
	.D5(output_8x10_o[4]),
	.D6(output_8x10_o[5]),
	.D7(output_8x10_o[6]),
	.D8(output_8x10_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x10_t_in),
	.TCE(1'd1),
	.OQ(output_8x10_pad_o),
	.TQ(output_8x10_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_14 (
	.I(output_8x10_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x10_t_out),
	.IO(dio1_p_6),
	.IOB(dio1_n_6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_60 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x11_o[0]),
	.D2(output_8x11_o[1]),
	.D3(output_8x11_o[2]),
	.D4(output_8x11_o[3]),
	.D5(output_8x11_o[4]),
	.D6(output_8x11_o[5]),
	.D7(output_8x11_o[6]),
	.D8(output_8x11_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x11_t_in),
	.TCE(1'd1),
	.OQ(output_8x11_pad_o),
	.TQ(output_8x11_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_15 (
	.I(output_8x11_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x11_t_out),
	.IO(dio1_p_7),
	.IOB(dio1_n_7)
);

OBUFTDS OBUFTDS_2(
	.I(spimaster0_interface_cs1[0]),
	.T(spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[0]),
	.OB(urukul2_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_3(
	.I(spimaster0_interface_cs1[1]),
	.T(spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[1]),
	.OB(urukul2_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_4(
	.I(spimaster0_interface_cs1[2]),
	.T(spimaster0_interface_offline),
	.O(urukul2_spi_p_cs_n[2]),
	.OB(urukul2_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_5(
	.I(spimaster0_interface_clk),
	.T(spimaster0_interface_offline),
	.O(urukul2_spi_p_clk),
	.OB(urukul2_spi_n_clk)
);

IOBUFDS IOBUFDS(
	.I(spimaster0_interface_sdo),
	.T((spimaster0_interface_offline | spimaster0_interface_half_duplex)),
	.IO(urukul2_spi_p_mosi),
	.IOB(urukul2_spi_n_mosi),
	.O(spimaster0_interface_mosi)
);

IOBUFDS IOBUFDS_1(
	.I(spimaster0_interface_sdo),
	.T(1'd1),
	.IO(urukul2_spi_p_miso),
	.IOB(urukul2_spi_n_miso),
	.O(spimaster0_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_61 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x12_o[0]),
	.D2(output_8x12_o[1]),
	.D3(output_8x12_o[2]),
	.D4(output_8x12_o[3]),
	.D5(output_8x12_o[4]),
	.D6(output_8x12_o[5]),
	.D7(output_8x12_o[6]),
	.D8(output_8x12_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x12_t_in),
	.TCE(1'd1),
	.OQ(output_8x12_pad_o),
	.TQ(output_8x12_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_16 (
	.I(output_8x12_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x12_t_out),
	.IO(urukul2_io_update_p),
	.IOB(urukul2_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_62 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x13_o[0]),
	.D2(output_8x13_o[1]),
	.D3(output_8x13_o[2]),
	.D4(output_8x13_o[3]),
	.D5(output_8x13_o[4]),
	.D6(output_8x13_o[5]),
	.D7(output_8x13_o[6]),
	.D8(output_8x13_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x13_t_in),
	.TCE(1'd1),
	.OQ(output_8x13_pad_o),
	.TQ(output_8x13_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_17 (
	.I(output_8x13_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x13_t_out),
	.IO(urukul2_sw0_p),
	.IOB(urukul2_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_63 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x14_o[0]),
	.D2(output_8x14_o[1]),
	.D3(output_8x14_o[2]),
	.D4(output_8x14_o[3]),
	.D5(output_8x14_o[4]),
	.D6(output_8x14_o[5]),
	.D7(output_8x14_o[6]),
	.D8(output_8x14_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x14_t_in),
	.TCE(1'd1),
	.OQ(output_8x14_pad_o),
	.TQ(output_8x14_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_18 (
	.I(output_8x14_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x14_t_out),
	.IO(urukul2_sw1_p),
	.IOB(urukul2_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_64 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x15_o[0]),
	.D2(output_8x15_o[1]),
	.D3(output_8x15_o[2]),
	.D4(output_8x15_o[3]),
	.D5(output_8x15_o[4]),
	.D6(output_8x15_o[5]),
	.D7(output_8x15_o[6]),
	.D8(output_8x15_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x15_t_in),
	.TCE(1'd1),
	.OQ(output_8x15_pad_o),
	.TQ(output_8x15_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_19 (
	.I(output_8x15_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x15_t_out),
	.IO(urukul2_sw2_p),
	.IOB(urukul2_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_65 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x16_o[0]),
	.D2(output_8x16_o[1]),
	.D3(output_8x16_o[2]),
	.D4(output_8x16_o[3]),
	.D5(output_8x16_o[4]),
	.D6(output_8x16_o[5]),
	.D7(output_8x16_o[6]),
	.D8(output_8x16_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x16_t_in),
	.TCE(1'd1),
	.OQ(output_8x16_pad_o),
	.TQ(output_8x16_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_20 (
	.I(output_8x16_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x16_t_out),
	.IO(urukul2_sw3_p),
	.IOB(urukul2_sw3_n)
);

OBUFTDS OBUFTDS_6(
	.I(spimaster1_interface_cs1[0]),
	.T(spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[0]),
	.OB(urukul4_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_7(
	.I(spimaster1_interface_cs1[1]),
	.T(spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[1]),
	.OB(urukul4_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_8(
	.I(spimaster1_interface_cs1[2]),
	.T(spimaster1_interface_offline),
	.O(urukul4_spi_p_cs_n[2]),
	.OB(urukul4_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_9(
	.I(spimaster1_interface_clk),
	.T(spimaster1_interface_offline),
	.O(urukul4_spi_p_clk),
	.OB(urukul4_spi_n_clk)
);

IOBUFDS IOBUFDS_2(
	.I(spimaster1_interface_sdo),
	.T((spimaster1_interface_offline | spimaster1_interface_half_duplex)),
	.IO(urukul4_spi_p_mosi),
	.IOB(urukul4_spi_n_mosi),
	.O(spimaster1_interface_mosi)
);

IOBUFDS IOBUFDS_3(
	.I(spimaster1_interface_sdo),
	.T(1'd1),
	.IO(urukul4_spi_p_miso),
	.IOB(urukul4_spi_n_miso),
	.O(spimaster1_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_66 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x17_o[0]),
	.D2(output_8x17_o[1]),
	.D3(output_8x17_o[2]),
	.D4(output_8x17_o[3]),
	.D5(output_8x17_o[4]),
	.D6(output_8x17_o[5]),
	.D7(output_8x17_o[6]),
	.D8(output_8x17_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x17_t_in),
	.TCE(1'd1),
	.OQ(output_8x17_pad_o),
	.TQ(output_8x17_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_21 (
	.I(output_8x17_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x17_t_out),
	.IO(urukul4_io_update_p),
	.IOB(urukul4_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_67 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x18_o[0]),
	.D2(output_8x18_o[1]),
	.D3(output_8x18_o[2]),
	.D4(output_8x18_o[3]),
	.D5(output_8x18_o[4]),
	.D6(output_8x18_o[5]),
	.D7(output_8x18_o[6]),
	.D8(output_8x18_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x18_t_in),
	.TCE(1'd1),
	.OQ(output_8x18_pad_o),
	.TQ(output_8x18_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_22 (
	.I(output_8x18_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x18_t_out),
	.IO(urukul4_sw0_p),
	.IOB(urukul4_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_68 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x19_o[0]),
	.D2(output_8x19_o[1]),
	.D3(output_8x19_o[2]),
	.D4(output_8x19_o[3]),
	.D5(output_8x19_o[4]),
	.D6(output_8x19_o[5]),
	.D7(output_8x19_o[6]),
	.D8(output_8x19_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x19_t_in),
	.TCE(1'd1),
	.OQ(output_8x19_pad_o),
	.TQ(output_8x19_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_23 (
	.I(output_8x19_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x19_t_out),
	.IO(urukul4_sw1_p),
	.IOB(urukul4_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_69 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x20_o[0]),
	.D2(output_8x20_o[1]),
	.D3(output_8x20_o[2]),
	.D4(output_8x20_o[3]),
	.D5(output_8x20_o[4]),
	.D6(output_8x20_o[5]),
	.D7(output_8x20_o[6]),
	.D8(output_8x20_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x20_t_in),
	.TCE(1'd1),
	.OQ(output_8x20_pad_o),
	.TQ(output_8x20_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_24 (
	.I(output_8x20_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x20_t_out),
	.IO(urukul4_sw2_p),
	.IOB(urukul4_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_70 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x21_o[0]),
	.D2(output_8x21_o[1]),
	.D3(output_8x21_o[2]),
	.D4(output_8x21_o[3]),
	.D5(output_8x21_o[4]),
	.D6(output_8x21_o[5]),
	.D7(output_8x21_o[6]),
	.D8(output_8x21_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x21_t_in),
	.TCE(1'd1),
	.OQ(output_8x21_pad_o),
	.TQ(output_8x21_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_25 (
	.I(output_8x21_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x21_t_out),
	.IO(urukul4_sw3_p),
	.IOB(urukul4_sw3_n)
);

OBUFTDS OBUFTDS_10(
	.I(spimaster2_interface_cs1[0]),
	.T(spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[0]),
	.OB(urukul6_spi_n_cs_n[0])
);

OBUFTDS OBUFTDS_11(
	.I(spimaster2_interface_cs1[1]),
	.T(spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[1]),
	.OB(urukul6_spi_n_cs_n[1])
);

OBUFTDS OBUFTDS_12(
	.I(spimaster2_interface_cs1[2]),
	.T(spimaster2_interface_offline),
	.O(urukul6_spi_p_cs_n[2]),
	.OB(urukul6_spi_n_cs_n[2])
);

OBUFTDS OBUFTDS_13(
	.I(spimaster2_interface_clk),
	.T(spimaster2_interface_offline),
	.O(urukul6_spi_p_clk),
	.OB(urukul6_spi_n_clk)
);

IOBUFDS IOBUFDS_4(
	.I(spimaster2_interface_sdo),
	.T((spimaster2_interface_offline | spimaster2_interface_half_duplex)),
	.IO(urukul6_spi_p_mosi),
	.IOB(urukul6_spi_n_mosi),
	.O(spimaster2_interface_mosi)
);

IOBUFDS IOBUFDS_5(
	.I(spimaster2_interface_sdo),
	.T(1'd1),
	.IO(urukul6_spi_p_miso),
	.IOB(urukul6_spi_n_miso),
	.O(spimaster2_interface_miso)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_71 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x22_o[0]),
	.D2(output_8x22_o[1]),
	.D3(output_8x22_o[2]),
	.D4(output_8x22_o[3]),
	.D5(output_8x22_o[4]),
	.D6(output_8x22_o[5]),
	.D7(output_8x22_o[6]),
	.D8(output_8x22_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x22_t_in),
	.TCE(1'd1),
	.OQ(output_8x22_pad_o),
	.TQ(output_8x22_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_26 (
	.I(output_8x22_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x22_t_out),
	.IO(urukul6_io_update_p),
	.IOB(urukul6_io_update_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_72 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x23_o[0]),
	.D2(output_8x23_o[1]),
	.D3(output_8x23_o[2]),
	.D4(output_8x23_o[3]),
	.D5(output_8x23_o[4]),
	.D6(output_8x23_o[5]),
	.D7(output_8x23_o[6]),
	.D8(output_8x23_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x23_t_in),
	.TCE(1'd1),
	.OQ(output_8x23_pad_o),
	.TQ(output_8x23_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_27 (
	.I(output_8x23_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x23_t_out),
	.IO(urukul6_sw0_p),
	.IOB(urukul6_sw0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_73 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x24_o[0]),
	.D2(output_8x24_o[1]),
	.D3(output_8x24_o[2]),
	.D4(output_8x24_o[3]),
	.D5(output_8x24_o[4]),
	.D6(output_8x24_o[5]),
	.D7(output_8x24_o[6]),
	.D8(output_8x24_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x24_t_in),
	.TCE(1'd1),
	.OQ(output_8x24_pad_o),
	.TQ(output_8x24_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_28 (
	.I(output_8x24_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x24_t_out),
	.IO(urukul6_sw1_p),
	.IOB(urukul6_sw1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_74 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x25_o[0]),
	.D2(output_8x25_o[1]),
	.D3(output_8x25_o[2]),
	.D4(output_8x25_o[3]),
	.D5(output_8x25_o[4]),
	.D6(output_8x25_o[5]),
	.D7(output_8x25_o[6]),
	.D8(output_8x25_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x25_t_in),
	.TCE(1'd1),
	.OQ(output_8x25_pad_o),
	.TQ(output_8x25_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_29 (
	.I(output_8x25_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x25_t_out),
	.IO(urukul6_sw2_p),
	.IOB(urukul6_sw2_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_75 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1(output_8x26_o[0]),
	.D2(output_8x26_o[1]),
	.D3(output_8x26_o[2]),
	.D4(output_8x26_o[3]),
	.D5(output_8x26_o[4]),
	.D6(output_8x26_o[5]),
	.D7(output_8x26_o[6]),
	.D8(output_8x26_o[7]),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(output_8x26_t_in),
	.TCE(1'd1),
	.OQ(output_8x26_pad_o),
	.TQ(output_8x26_t_out)
);

IOBUFDS_INTERMDISABLE #(
	.DIFF_TERM("FALSE"),
	.IBUF_LOW_PWR("TRUE"),
	.USE_IBUFDISABLE("TRUE")
) IOBUFDS_INTERMDISABLE_30 (
	.I(output_8x26_pad_o),
	.IBUFDISABLE(1'd1),
	.INTERMDISABLE(1'd1),
	.T(output_8x26_t_out),
	.IO(urukul6_sw3_p),
	.IOB(urukul6_sw3_n)
);

IBUFGDS #(
	.DIFF_TERM("TRUE"),
	.IBUF_LOW_PWR("FALSE")
) IBUFGDS (
	.I(si5324_clkout_fabric_p),
	.IB(si5324_clkout_fabric_n),
	.O(monroe_ionphoton_rtio_crg_clk_synth_se)
);

PLLE2_ADV #(
	.BANDWIDTH("HIGH"),
	.CLKFBOUT_MULT(4'd12),
	.CLKIN1_PERIOD(8.0),
	.CLKIN2_PERIOD(8.0),
	.CLKOUT0_DIVIDE(2'd3),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd12),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.001),
	.STARTUP_WAIT("FALSE")
) PLLE2_ADV (
	.CLKFBIN(monroe_ionphoton_rtio_crg_fb_clk),
	.CLKIN2(monroe_ionphoton_rtio_crg_clk_synth_se),
	.CLKINSEL(1'd0),
	.RST(monroe_ionphoton_rtio_crg_storage),
	.CLKFBOUT(monroe_ionphoton_rtio_crg_fb_clk),
	.CLKOUT0(monroe_ionphoton_rtio_crg_rtiox4_clk),
	.CLKOUT1(monroe_ionphoton_rtio_crg_rtio_clk),
	.LOCKED(monroe_ionphoton_rtio_crg_pll_locked)
);

BUFG BUFG_8(
	.I(monroe_ionphoton_rtio_crg_rtio_clk),
	.O(rtio_clk)
);

BUFG BUFG_9(
	.I(monroe_ionphoton_rtio_crg_rtiox4_clk),
	.O(rtiox4_clk)
);

reg [13:0] latency_compensation[0:36];
reg [5:0] memadr_15;
always @(posedge rsys_clk) begin
	memadr_15 <= monroe_ionphoton_rtio_core_outputs_lanedistributor_adr;
end

assign monroe_ionphoton_rtio_core_outputs_lanedistributor_dat_r = latency_compensation[memadr_15];

initial begin
	$readmemh("latency_compensation.init", latency_compensation);
end

reg [115:0] storage_7[0:127];
reg [6:0] memadr_16;
reg [6:0] memadr_17;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_we)
		storage_7[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
	memadr_16 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_17 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r = storage_7[memadr_16];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r = storage_7[memadr_17];

reg [115:0] storage_8[0:127];
reg [6:0] memadr_18;
reg [6:0] memadr_19;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_we)
		storage_8[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
	memadr_18 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_19 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r = storage_8[memadr_18];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r = storage_8[memadr_19];

reg [115:0] storage_9[0:127];
reg [6:0] memadr_20;
reg [6:0] memadr_21;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_we)
		storage_9[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
	memadr_20 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_21 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r = storage_9[memadr_20];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r = storage_9[memadr_21];

reg [115:0] storage_10[0:127];
reg [6:0] memadr_22;
reg [6:0] memadr_23;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_we)
		storage_10[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
	memadr_22 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_23 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r = storage_10[memadr_22];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r = storage_10[memadr_23];

reg [115:0] storage_11[0:127];
reg [6:0] memadr_24;
reg [6:0] memadr_25;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_we)
		storage_11[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
	memadr_24 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_25 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r = storage_11[memadr_24];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r = storage_11[memadr_25];

reg [115:0] storage_12[0:127];
reg [6:0] memadr_26;
reg [6:0] memadr_27;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_we)
		storage_12[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
	memadr_26 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_27 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r = storage_12[memadr_26];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r = storage_12[memadr_27];

reg [115:0] storage_13[0:127];
reg [6:0] memadr_28;
reg [6:0] memadr_29;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_we)
		storage_13[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
	memadr_28 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_29 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r = storage_13[memadr_28];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r = storage_13[memadr_29];

reg [115:0] storage_14[0:127];
reg [6:0] memadr_30;
reg [6:0] memadr_31;
always @(posedge rsys_clk) begin
	if (monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_we)
		storage_14[monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_adr] <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
	memadr_30 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_31 <= monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
end

assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r = storage_14[memadr_30];
assign monroe_ionphoton_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r = storage_14[memadr_31];

reg [0:0] en_replaces_rom[0:36];
reg [5:0] memadr_32;
always @(posedge rio_clk) begin
	memadr_32 <= monroe_ionphoton_rtio_core_outputs_memory0_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory0_dat_r = en_replaces_rom[memadr_32];

initial begin
	$readmemh("en_replaces_rom.init", en_replaces_rom);
end

reg [0:0] en_replaces_rom_1[0:36];
reg [5:0] memadr_33;
always @(posedge rio_clk) begin
	memadr_33 <= monroe_ionphoton_rtio_core_outputs_memory1_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory1_dat_r = en_replaces_rom_1[memadr_33];

initial begin
	$readmemh("en_replaces_rom_1.init", en_replaces_rom_1);
end

reg [0:0] en_replaces_rom_2[0:36];
reg [5:0] memadr_34;
always @(posedge rio_clk) begin
	memadr_34 <= monroe_ionphoton_rtio_core_outputs_memory2_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory2_dat_r = en_replaces_rom_2[memadr_34];

initial begin
	$readmemh("en_replaces_rom_2.init", en_replaces_rom_2);
end

reg [0:0] en_replaces_rom_3[0:36];
reg [5:0] memadr_35;
always @(posedge rio_clk) begin
	memadr_35 <= monroe_ionphoton_rtio_core_outputs_memory3_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory3_dat_r = en_replaces_rom_3[memadr_35];

initial begin
	$readmemh("en_replaces_rom_3.init", en_replaces_rom_3);
end

reg [0:0] en_replaces_rom_4[0:36];
reg [5:0] memadr_36;
always @(posedge rio_clk) begin
	memadr_36 <= monroe_ionphoton_rtio_core_outputs_memory4_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory4_dat_r = en_replaces_rom_4[memadr_36];

initial begin
	$readmemh("en_replaces_rom_4.init", en_replaces_rom_4);
end

reg [0:0] en_replaces_rom_5[0:36];
reg [5:0] memadr_37;
always @(posedge rio_clk) begin
	memadr_37 <= monroe_ionphoton_rtio_core_outputs_memory5_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory5_dat_r = en_replaces_rom_5[memadr_37];

initial begin
	$readmemh("en_replaces_rom_5.init", en_replaces_rom_5);
end

reg [0:0] en_replaces_rom_6[0:36];
reg [5:0] memadr_38;
always @(posedge rio_clk) begin
	memadr_38 <= monroe_ionphoton_rtio_core_outputs_memory6_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory6_dat_r = en_replaces_rom_6[memadr_38];

initial begin
	$readmemh("en_replaces_rom_6.init", en_replaces_rom_6);
end

reg [0:0] en_replaces_rom_7[0:36];
reg [5:0] memadr_39;
always @(posedge rio_clk) begin
	memadr_39 <= monroe_ionphoton_rtio_core_outputs_memory7_adr;
end

assign monroe_ionphoton_rtio_core_outputs_memory7_dat_r = en_replaces_rom_7[memadr_39];

initial begin
	$readmemh("en_replaces_rom_7.init", en_replaces_rom_7);
end

reg [64:0] storage_15[0:63];
reg [5:0] memadr_40;
reg [5:0] memadr_41;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_we)
		storage_15[monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_dat_w;
	memadr_40 <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_41 <= monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_wrport_dat_r = storage_15[memadr_40];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo0_rdport_dat_r = storage_15[memadr_41];

reg [64:0] storage_16[0:63];
reg [5:0] memadr_42;
reg [5:0] memadr_43;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_we)
		storage_16[monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_dat_w;
	memadr_42 <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_43 <= monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_wrport_dat_r = storage_16[memadr_42];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo1_rdport_dat_r = storage_16[memadr_43];

reg [64:0] storage_17[0:63];
reg [5:0] memadr_44;
reg [5:0] memadr_45;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_we)
		storage_17[monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_dat_w;
	memadr_44 <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_45 <= monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_wrport_dat_r = storage_17[memadr_44];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo2_rdport_dat_r = storage_17[memadr_45];

reg [64:0] storage_18[0:63];
reg [5:0] memadr_46;
reg [5:0] memadr_47;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_we)
		storage_18[monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_dat_w;
	memadr_46 <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_47 <= monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_wrport_dat_r = storage_18[memadr_46];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo3_rdport_dat_r = storage_18[memadr_47];

reg [31:0] storage_19[0:3];
reg [1:0] memadr_48;
reg [1:0] memadr_49;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_we)
		storage_19[monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_dat_w;
	memadr_48 <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_49 <= monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_wrport_dat_r = storage_19[memadr_48];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo4_rdport_dat_r = storage_19[memadr_49];

reg [31:0] storage_20[0:3];
reg [1:0] memadr_50;
reg [1:0] memadr_51;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_we)
		storage_20[monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_dat_w;
	memadr_50 <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_51 <= monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_wrport_dat_r = storage_20[memadr_50];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo5_rdport_dat_r = storage_20[memadr_51];

reg [31:0] storage_21[0:3];
reg [1:0] memadr_52;
reg [1:0] memadr_53;
always @(posedge rio_clk) begin
	if (monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_we)
		storage_21[monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_adr] <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_dat_w;
	memadr_52 <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_53 <= monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_adr;
end

assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_wrport_dat_r = storage_21[memadr_52];
assign monroe_ionphoton_rtio_core_inputs_asyncfifo6_rdport_dat_r = storage_21[memadr_53];

reg [256:0] storage_22[0:127];
reg [256:0] memdat_5;
reg [256:0] memdat_6;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_rtio_analyzer_fifo_wrport_we)
		storage_22[monroe_ionphoton_rtio_analyzer_fifo_wrport_adr] <= monroe_ionphoton_rtio_analyzer_fifo_wrport_dat_w;
	memdat_5 <= storage_22[monroe_ionphoton_rtio_analyzer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_rtio_analyzer_fifo_rdport_re)
		memdat_6 <= storage_22[monroe_ionphoton_rtio_analyzer_fifo_rdport_adr];
end

assign monroe_ionphoton_rtio_analyzer_fifo_wrport_dat_r = memdat_5;
assign monroe_ionphoton_rtio_analyzer_fifo_rdport_dat_r = memdat_6;

reg [7:0] data_mem_grain0[0:8191];
reg [12:0] memadr_54;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[0])
		data_mem_grain0[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[7:0];
	memadr_54 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[7:0] = data_mem_grain0[memadr_54];

reg [7:0] data_mem_grain1[0:8191];
reg [12:0] memadr_55;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[1])
		data_mem_grain1[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[15:8];
	memadr_55 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[15:8] = data_mem_grain1[memadr_55];

reg [7:0] data_mem_grain2[0:8191];
reg [12:0] memadr_56;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[2])
		data_mem_grain2[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[23:16];
	memadr_56 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[23:16] = data_mem_grain2[memadr_56];

reg [7:0] data_mem_grain3[0:8191];
reg [12:0] memadr_57;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[3])
		data_mem_grain3[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[31:24];
	memadr_57 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[31:24] = data_mem_grain3[memadr_57];

reg [7:0] data_mem_grain4[0:8191];
reg [12:0] memadr_58;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[4])
		data_mem_grain4[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[39:32];
	memadr_58 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[39:32] = data_mem_grain4[memadr_58];

reg [7:0] data_mem_grain5[0:8191];
reg [12:0] memadr_59;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[5])
		data_mem_grain5[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[47:40];
	memadr_59 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[47:40] = data_mem_grain5[memadr_59];

reg [7:0] data_mem_grain6[0:8191];
reg [12:0] memadr_60;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[6])
		data_mem_grain6[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[55:48];
	memadr_60 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[55:48] = data_mem_grain6[memadr_60];

reg [7:0] data_mem_grain7[0:8191];
reg [12:0] memadr_61;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[7])
		data_mem_grain7[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[63:56];
	memadr_61 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[63:56] = data_mem_grain7[memadr_61];

reg [7:0] data_mem_grain8[0:8191];
reg [12:0] memadr_62;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[8])
		data_mem_grain8[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[71:64];
	memadr_62 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[71:64] = data_mem_grain8[memadr_62];

reg [7:0] data_mem_grain9[0:8191];
reg [12:0] memadr_63;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[9])
		data_mem_grain9[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[79:72];
	memadr_63 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[79:72] = data_mem_grain9[memadr_63];

reg [7:0] data_mem_grain10[0:8191];
reg [12:0] memadr_64;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[10])
		data_mem_grain10[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[87:80];
	memadr_64 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[87:80] = data_mem_grain10[memadr_64];

reg [7:0] data_mem_grain11[0:8191];
reg [12:0] memadr_65;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[11])
		data_mem_grain11[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[95:88];
	memadr_65 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[95:88] = data_mem_grain11[memadr_65];

reg [7:0] data_mem_grain12[0:8191];
reg [12:0] memadr_66;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[12])
		data_mem_grain12[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[103:96];
	memadr_66 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[103:96] = data_mem_grain12[memadr_66];

reg [7:0] data_mem_grain13[0:8191];
reg [12:0] memadr_67;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[13])
		data_mem_grain13[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[111:104];
	memadr_67 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[111:104] = data_mem_grain13[memadr_67];

reg [7:0] data_mem_grain14[0:8191];
reg [12:0] memadr_68;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[14])
		data_mem_grain14[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[119:112];
	memadr_68 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[119:112] = data_mem_grain14[memadr_68];

reg [7:0] data_mem_grain15[0:8191];
reg [12:0] memadr_69;
always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_we[15])
		data_mem_grain15[monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr] <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_w[127:120];
	memadr_69 <= monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_adr;
end

assign monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_monroe_ionphoton_data_port_dat_r[127:120] = data_mem_grain15[memadr_69];

reg [7:0] mem_grain0[0:381];
reg [8:0] memadr_70;
reg [8:0] memadr_71;
always @(posedge sys_clk) begin
	memadr_70 <= monroe_ionphoton_monroe_ionphoton_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram0_we[0])
		mem_grain0[monroe_ionphoton_monroe_ionphoton_sram0_adr1] <= monroe_ionphoton_monroe_ionphoton_sram0_dat_w[7:0];
	memadr_71 <= monroe_ionphoton_monroe_ionphoton_sram0_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r[7:0] = mem_grain0[memadr_70];
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_r1[7:0] = mem_grain0[memadr_71];

reg [7:0] mem_grain1[0:381];
reg [8:0] memadr_72;
reg [8:0] memadr_73;
always @(posedge sys_clk) begin
	memadr_72 <= monroe_ionphoton_monroe_ionphoton_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram0_we[1])
		mem_grain1[monroe_ionphoton_monroe_ionphoton_sram0_adr1] <= monroe_ionphoton_monroe_ionphoton_sram0_dat_w[15:8];
	memadr_73 <= monroe_ionphoton_monroe_ionphoton_sram0_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r[15:8] = mem_grain1[memadr_72];
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_r1[15:8] = mem_grain1[memadr_73];

reg [7:0] mem_grain2[0:381];
reg [8:0] memadr_74;
reg [8:0] memadr_75;
always @(posedge sys_clk) begin
	memadr_74 <= monroe_ionphoton_monroe_ionphoton_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram0_we[2])
		mem_grain2[monroe_ionphoton_monroe_ionphoton_sram0_adr1] <= monroe_ionphoton_monroe_ionphoton_sram0_dat_w[23:16];
	memadr_75 <= monroe_ionphoton_monroe_ionphoton_sram0_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r[23:16] = mem_grain2[memadr_74];
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_r1[23:16] = mem_grain2[memadr_75];

reg [7:0] mem_grain3[0:381];
reg [8:0] memadr_76;
reg [8:0] memadr_77;
always @(posedge sys_clk) begin
	memadr_76 <= monroe_ionphoton_monroe_ionphoton_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram0_we[3])
		mem_grain3[monroe_ionphoton_monroe_ionphoton_sram0_adr1] <= monroe_ionphoton_monroe_ionphoton_sram0_dat_w[31:24];
	memadr_77 <= monroe_ionphoton_monroe_ionphoton_sram0_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory0_dat_r[31:24] = mem_grain3[memadr_76];
assign monroe_ionphoton_monroe_ionphoton_sram0_dat_r1[31:24] = mem_grain3[memadr_77];

reg [7:0] mem_grain0_1[0:381];
reg [8:0] memadr_78;
reg [8:0] memadr_79;
always @(posedge sys_clk) begin
	memadr_78 <= monroe_ionphoton_monroe_ionphoton_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram1_we[0])
		mem_grain0_1[monroe_ionphoton_monroe_ionphoton_sram1_adr1] <= monroe_ionphoton_monroe_ionphoton_sram1_dat_w[7:0];
	memadr_79 <= monroe_ionphoton_monroe_ionphoton_sram1_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r[7:0] = mem_grain0_1[memadr_78];
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_r1[7:0] = mem_grain0_1[memadr_79];

reg [7:0] mem_grain1_1[0:381];
reg [8:0] memadr_80;
reg [8:0] memadr_81;
always @(posedge sys_clk) begin
	memadr_80 <= monroe_ionphoton_monroe_ionphoton_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram1_we[1])
		mem_grain1_1[monroe_ionphoton_monroe_ionphoton_sram1_adr1] <= monroe_ionphoton_monroe_ionphoton_sram1_dat_w[15:8];
	memadr_81 <= monroe_ionphoton_monroe_ionphoton_sram1_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r[15:8] = mem_grain1_1[memadr_80];
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_r1[15:8] = mem_grain1_1[memadr_81];

reg [7:0] mem_grain2_1[0:381];
reg [8:0] memadr_82;
reg [8:0] memadr_83;
always @(posedge sys_clk) begin
	memadr_82 <= monroe_ionphoton_monroe_ionphoton_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram1_we[2])
		mem_grain2_1[monroe_ionphoton_monroe_ionphoton_sram1_adr1] <= monroe_ionphoton_monroe_ionphoton_sram1_dat_w[23:16];
	memadr_83 <= monroe_ionphoton_monroe_ionphoton_sram1_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r[23:16] = mem_grain2_1[memadr_82];
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_r1[23:16] = mem_grain2_1[memadr_83];

reg [7:0] mem_grain3_1[0:381];
reg [8:0] memadr_84;
reg [8:0] memadr_85;
always @(posedge sys_clk) begin
	memadr_84 <= monroe_ionphoton_monroe_ionphoton_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram1_we[3])
		mem_grain3_1[monroe_ionphoton_monroe_ionphoton_sram1_adr1] <= monroe_ionphoton_monroe_ionphoton_sram1_dat_w[31:24];
	memadr_85 <= monroe_ionphoton_monroe_ionphoton_sram1_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory1_dat_r[31:24] = mem_grain3_1[memadr_84];
assign monroe_ionphoton_monroe_ionphoton_sram1_dat_r1[31:24] = mem_grain3_1[memadr_85];

reg [7:0] mem_grain0_2[0:381];
reg [8:0] memadr_86;
reg [8:0] memadr_87;
always @(posedge sys_clk) begin
	memadr_86 <= monroe_ionphoton_monroe_ionphoton_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram2_we[0])
		mem_grain0_2[monroe_ionphoton_monroe_ionphoton_sram2_adr1] <= monroe_ionphoton_monroe_ionphoton_sram2_dat_w[7:0];
	memadr_87 <= monroe_ionphoton_monroe_ionphoton_sram2_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r[7:0] = mem_grain0_2[memadr_86];
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_r1[7:0] = mem_grain0_2[memadr_87];

reg [7:0] mem_grain1_2[0:381];
reg [8:0] memadr_88;
reg [8:0] memadr_89;
always @(posedge sys_clk) begin
	memadr_88 <= monroe_ionphoton_monroe_ionphoton_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram2_we[1])
		mem_grain1_2[monroe_ionphoton_monroe_ionphoton_sram2_adr1] <= monroe_ionphoton_monroe_ionphoton_sram2_dat_w[15:8];
	memadr_89 <= monroe_ionphoton_monroe_ionphoton_sram2_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r[15:8] = mem_grain1_2[memadr_88];
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_r1[15:8] = mem_grain1_2[memadr_89];

reg [7:0] mem_grain2_2[0:381];
reg [8:0] memadr_90;
reg [8:0] memadr_91;
always @(posedge sys_clk) begin
	memadr_90 <= monroe_ionphoton_monroe_ionphoton_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram2_we[2])
		mem_grain2_2[monroe_ionphoton_monroe_ionphoton_sram2_adr1] <= monroe_ionphoton_monroe_ionphoton_sram2_dat_w[23:16];
	memadr_91 <= monroe_ionphoton_monroe_ionphoton_sram2_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r[23:16] = mem_grain2_2[memadr_90];
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_r1[23:16] = mem_grain2_2[memadr_91];

reg [7:0] mem_grain3_2[0:381];
reg [8:0] memadr_92;
reg [8:0] memadr_93;
always @(posedge sys_clk) begin
	memadr_92 <= monroe_ionphoton_monroe_ionphoton_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram2_we[3])
		mem_grain3_2[monroe_ionphoton_monroe_ionphoton_sram2_adr1] <= monroe_ionphoton_monroe_ionphoton_sram2_dat_w[31:24];
	memadr_93 <= monroe_ionphoton_monroe_ionphoton_sram2_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory2_dat_r[31:24] = mem_grain3_2[memadr_92];
assign monroe_ionphoton_monroe_ionphoton_sram2_dat_r1[31:24] = mem_grain3_2[memadr_93];

reg [7:0] mem_grain0_3[0:381];
reg [8:0] memadr_94;
reg [8:0] memadr_95;
always @(posedge sys_clk) begin
	memadr_94 <= monroe_ionphoton_monroe_ionphoton_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram3_we[0])
		mem_grain0_3[monroe_ionphoton_monroe_ionphoton_sram3_adr1] <= monroe_ionphoton_monroe_ionphoton_sram3_dat_w[7:0];
	memadr_95 <= monroe_ionphoton_monroe_ionphoton_sram3_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r[7:0] = mem_grain0_3[memadr_94];
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_r1[7:0] = mem_grain0_3[memadr_95];

reg [7:0] mem_grain1_3[0:381];
reg [8:0] memadr_96;
reg [8:0] memadr_97;
always @(posedge sys_clk) begin
	memadr_96 <= monroe_ionphoton_monroe_ionphoton_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram3_we[1])
		mem_grain1_3[monroe_ionphoton_monroe_ionphoton_sram3_adr1] <= monroe_ionphoton_monroe_ionphoton_sram3_dat_w[15:8];
	memadr_97 <= monroe_ionphoton_monroe_ionphoton_sram3_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r[15:8] = mem_grain1_3[memadr_96];
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_r1[15:8] = mem_grain1_3[memadr_97];

reg [7:0] mem_grain2_3[0:381];
reg [8:0] memadr_98;
reg [8:0] memadr_99;
always @(posedge sys_clk) begin
	memadr_98 <= monroe_ionphoton_monroe_ionphoton_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram3_we[2])
		mem_grain2_3[monroe_ionphoton_monroe_ionphoton_sram3_adr1] <= monroe_ionphoton_monroe_ionphoton_sram3_dat_w[23:16];
	memadr_99 <= monroe_ionphoton_monroe_ionphoton_sram3_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r[23:16] = mem_grain2_3[memadr_98];
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_r1[23:16] = mem_grain2_3[memadr_99];

reg [7:0] mem_grain3_3[0:381];
reg [8:0] memadr_100;
reg [8:0] memadr_101;
always @(posedge sys_clk) begin
	memadr_100 <= monroe_ionphoton_monroe_ionphoton_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (monroe_ionphoton_monroe_ionphoton_sram3_we[3])
		mem_grain3_3[monroe_ionphoton_monroe_ionphoton_sram3_adr1] <= monroe_ionphoton_monroe_ionphoton_sram3_dat_w[31:24];
	memadr_101 <= monroe_ionphoton_monroe_ionphoton_sram3_adr1;
end

assign monroe_ionphoton_monroe_ionphoton_reader_memory3_dat_r[31:24] = mem_grain3_3[memadr_100];
assign monroe_ionphoton_monroe_ionphoton_sram3_dat_r1[31:24] = mem_grain3_3[memadr_101];

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(clk200_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(eth_tx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(eth_rx_rst)
);

OBUFDS OBUFDS_1(
	.I(pad0),
	.O(urukul2_dds_reset_sync_in_p),
	.OB(urukul2_dds_reset_sync_in_n)
);

OBUFDS OBUFDS_2(
	.I(pad1),
	.O(urukul4_dds_reset_sync_in_p),
	.OB(urukul4_dds_reset_sync_in_n)
);

OBUFDS OBUFDS_3(
	.I(pad2),
	.O(urukul6_dds_reset_sync_in_p),
	.OB(urukul6_dds_reset_sync_in_n)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl3),
	.Q(xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl3),
	.Q(rtio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(rio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(monroe_ionphoton_rtio_core_cmd_reset),
	.Q(xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(rio_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(monroe_ionphoton_rtio_core_cmd_reset),
	.Q(rio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(monroe_ionphoton_rtio_core_cmd_reset_phy),
	.Q(xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(monroe_ionphoton_rtio_core_cmd_reset_phy),
	.Q(rio_phy_rst)
);

endmodule
